// Created by ihdl
module Data_Bank ( clk, write, dira, data, A, dirb, B );
  input [4:0] dira;
  input [23:0] data;
  output [23:0] A;
  input [4:0] dirb;
  output [23:0] B;
  input clk, write;
  wire   \mem[0][23] , \mem[0][22] , \mem[0][21] , \mem[0][20] , \mem[0][19] ,
         \mem[0][18] , \mem[0][17] , \mem[0][16] , \mem[0][15] , \mem[0][14] ,
         \mem[0][13] , \mem[0][12] , \mem[0][11] , \mem[0][10] , \mem[0][9] ,
         \mem[0][8] , \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] ,
         \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , \mem[1][23] ,
         \mem[1][22] , \mem[1][21] , \mem[1][20] , \mem[1][19] , \mem[1][18] ,
         \mem[1][17] , \mem[1][16] , \mem[1][15] , \mem[1][14] , \mem[1][13] ,
         \mem[1][12] , \mem[1][11] , \mem[1][10] , \mem[1][9] , \mem[1][8] ,
         \mem[1][7] , \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] ,
         \mem[1][2] , \mem[1][1] , \mem[1][0] , \mem[2][23] , \mem[2][22] ,
         \mem[2][21] , \mem[2][20] , \mem[2][19] , \mem[2][18] , \mem[2][17] ,
         \mem[2][16] , \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] ,
         \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[3][23] , \mem[3][22] , \mem[3][21] ,
         \mem[3][20] , \mem[3][19] , \mem[3][18] , \mem[3][17] , \mem[3][16] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[4][23] , \mem[4][22] , \mem[4][21] , \mem[4][20] ,
         \mem[4][19] , \mem[4][18] , \mem[4][17] , \mem[4][16] , \mem[4][15] ,
         \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] , \mem[4][10] ,
         \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] , \mem[4][5] ,
         \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] , \mem[4][0] ,
         \mem[5][23] , \mem[5][22] , \mem[5][21] , \mem[5][20] , \mem[5][19] ,
         \mem[5][18] , \mem[5][17] , \mem[5][16] , \mem[5][15] , \mem[5][14] ,
         \mem[5][13] , \mem[5][12] , \mem[5][11] , \mem[5][10] , \mem[5][9] ,
         \mem[5][8] , \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] ,
         \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[6][23] ,
         \mem[6][22] , \mem[6][21] , \mem[6][20] , \mem[6][19] , \mem[6][18] ,
         \mem[6][17] , \mem[6][16] , \mem[6][15] , \mem[6][14] , \mem[6][13] ,
         \mem[6][12] , \mem[6][11] , \mem[6][10] , \mem[6][9] , \mem[6][8] ,
         \mem[6][7] , \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] ,
         \mem[6][2] , \mem[6][1] , \mem[6][0] , \mem[7][23] , \mem[7][22] ,
         \mem[7][21] , \mem[7][20] , \mem[7][19] , \mem[7][18] , \mem[7][17] ,
         \mem[7][16] , \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] ,
         \mem[7][11] , \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[8][23] , \mem[8][22] , \mem[8][21] ,
         \mem[8][20] , \mem[8][19] , \mem[8][18] , \mem[8][17] , \mem[8][16] ,
         \mem[8][15] , \mem[8][14] , \mem[8][13] , \mem[8][12] , \mem[8][11] ,
         \mem[8][10] , \mem[8][9] , \mem[8][8] , \mem[8][7] , \mem[8][6] ,
         \mem[8][5] , \mem[8][4] , \mem[8][3] , \mem[8][2] , \mem[8][1] ,
         \mem[8][0] , \mem[9][23] , \mem[9][22] , \mem[9][21] , \mem[9][20] ,
         \mem[9][19] , \mem[9][18] , \mem[9][17] , \mem[9][16] , \mem[9][15] ,
         \mem[9][14] , \mem[9][13] , \mem[9][12] , \mem[9][11] , \mem[9][10] ,
         \mem[9][9] , \mem[9][8] , \mem[9][7] , \mem[9][6] , \mem[9][5] ,
         \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] , \mem[9][0] ,
         \mem[10][23] , \mem[10][22] , \mem[10][21] , \mem[10][20] ,
         \mem[10][19] , \mem[10][18] , \mem[10][17] , \mem[10][16] ,
         \mem[10][15] , \mem[10][14] , \mem[10][13] , \mem[10][12] ,
         \mem[10][11] , \mem[10][10] , \mem[10][9] , \mem[10][8] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[11][23] ,
         \mem[11][22] , \mem[11][21] , \mem[11][20] , \mem[11][19] ,
         \mem[11][18] , \mem[11][17] , \mem[11][16] , \mem[11][15] ,
         \mem[11][14] , \mem[11][13] , \mem[11][12] , \mem[11][11] ,
         \mem[11][10] , \mem[11][9] , \mem[11][8] , \mem[11][7] , \mem[11][6] ,
         \mem[11][5] , \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] ,
         \mem[11][0] , \mem[12][23] , \mem[12][22] , \mem[12][21] ,
         \mem[12][20] , \mem[12][19] , \mem[12][18] , \mem[12][17] ,
         \mem[12][16] , \mem[12][15] , \mem[12][14] , \mem[12][13] ,
         \mem[12][12] , \mem[12][11] , \mem[12][10] , \mem[12][9] ,
         \mem[12][8] , \mem[12][7] , \mem[12][6] , \mem[12][5] , \mem[12][4] ,
         \mem[12][3] , \mem[12][2] , \mem[12][1] , \mem[12][0] , \mem[13][23] ,
         \mem[13][22] , \mem[13][21] , \mem[13][20] , \mem[13][19] ,
         \mem[13][18] , \mem[13][17] , \mem[13][16] , \mem[13][15] ,
         \mem[13][14] , \mem[13][13] , \mem[13][12] , \mem[13][11] ,
         \mem[13][10] , \mem[13][9] , \mem[13][8] , \mem[13][7] , \mem[13][6] ,
         \mem[13][5] , \mem[13][4] , \mem[13][3] , \mem[13][2] , \mem[13][1] ,
         \mem[13][0] , \mem[14][23] , \mem[14][22] , \mem[14][21] ,
         \mem[14][20] , \mem[14][19] , \mem[14][18] , \mem[14][17] ,
         \mem[14][16] , \mem[14][15] , \mem[14][14] , \mem[14][13] ,
         \mem[14][12] , \mem[14][11] , \mem[14][10] , \mem[14][9] ,
         \mem[14][8] , \mem[14][7] , \mem[14][6] , \mem[14][5] , \mem[14][4] ,
         \mem[14][3] , \mem[14][2] , \mem[14][1] , \mem[14][0] , \mem[15][23] ,
         \mem[15][22] , \mem[15][21] , \mem[15][20] , \mem[15][19] ,
         \mem[15][18] , \mem[15][17] , \mem[15][16] , \mem[15][15] ,
         \mem[15][14] , \mem[15][13] , \mem[15][12] , \mem[15][11] ,
         \mem[15][10] , \mem[15][9] , \mem[15][8] , \mem[15][7] , \mem[15][6] ,
         \mem[15][5] , \mem[15][4] , \mem[15][3] , \mem[15][2] , \mem[15][1] ,
         \mem[15][0] , \mem[16][23] , \mem[16][22] , \mem[16][21] ,
         \mem[16][20] , \mem[16][19] , \mem[16][18] , \mem[16][17] ,
         \mem[16][16] , \mem[16][15] , \mem[16][14] , \mem[16][13] ,
         \mem[16][12] , \mem[16][11] , \mem[16][10] , \mem[16][9] ,
         \mem[16][8] , \mem[16][7] , \mem[16][6] , \mem[16][5] , \mem[16][4] ,
         \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] , \mem[17][23] ,
         \mem[17][22] , \mem[17][21] , \mem[17][20] , \mem[17][19] ,
         \mem[17][18] , \mem[17][17] , \mem[17][16] , \mem[17][15] ,
         \mem[17][14] , \mem[17][13] , \mem[17][12] , \mem[17][11] ,
         \mem[17][10] , \mem[17][9] , \mem[17][8] , \mem[17][7] , \mem[17][6] ,
         \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] , \mem[17][1] ,
         \mem[17][0] , \mem[18][23] , \mem[18][22] , \mem[18][21] ,
         \mem[18][20] , \mem[18][19] , \mem[18][18] , \mem[18][17] ,
         \mem[18][16] , \mem[18][15] , \mem[18][14] , \mem[18][13] ,
         \mem[18][12] , \mem[18][11] , \mem[18][10] , \mem[18][9] ,
         \mem[18][8] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[19][23] ,
         \mem[19][22] , \mem[19][21] , \mem[19][20] , \mem[19][19] ,
         \mem[19][18] , \mem[19][17] , \mem[19][16] , \mem[19][15] ,
         \mem[19][14] , \mem[19][13] , \mem[19][12] , \mem[19][11] ,
         \mem[19][10] , \mem[19][9] , \mem[19][8] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[20][23] , \mem[20][22] , \mem[20][21] ,
         \mem[20][20] , \mem[20][19] , \mem[20][18] , \mem[20][17] ,
         \mem[20][16] , \mem[20][15] , \mem[20][14] , \mem[20][13] ,
         \mem[20][12] , \mem[20][11] , \mem[20][10] , \mem[20][9] ,
         \mem[20][8] , \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] ,
         \mem[20][3] , \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[21][23] ,
         \mem[21][22] , \mem[21][21] , \mem[21][20] , \mem[21][19] ,
         \mem[21][18] , \mem[21][17] , \mem[21][16] , \mem[21][15] ,
         \mem[21][14] , \mem[21][13] , \mem[21][12] , \mem[21][11] ,
         \mem[21][10] , \mem[21][9] , \mem[21][8] , \mem[21][7] , \mem[21][6] ,
         \mem[21][5] , \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] ,
         \mem[21][0] , \mem[22][23] , \mem[22][22] , \mem[22][21] ,
         \mem[22][20] , \mem[22][19] , \mem[22][18] , \mem[22][17] ,
         \mem[22][16] , \mem[22][15] , \mem[22][14] , \mem[22][13] ,
         \mem[22][12] , \mem[22][11] , \mem[22][10] , \mem[22][9] ,
         \mem[22][8] , \mem[22][7] , \mem[22][6] , \mem[22][5] , \mem[22][4] ,
         \mem[22][3] , \mem[22][2] , \mem[22][1] , \mem[22][0] , \mem[23][23] ,
         \mem[23][22] , \mem[23][21] , \mem[23][20] , \mem[23][19] ,
         \mem[23][18] , \mem[23][17] , \mem[23][16] , \mem[23][15] ,
         \mem[23][14] , \mem[23][13] , \mem[23][12] , \mem[23][11] ,
         \mem[23][10] , \mem[23][9] , \mem[23][8] , \mem[23][7] , \mem[23][6] ,
         \mem[23][5] , \mem[23][4] , \mem[23][3] , \mem[23][2] , \mem[23][1] ,
         \mem[23][0] , \mem[24][23] , \mem[24][22] , \mem[24][21] ,
         \mem[24][20] , \mem[24][19] , \mem[24][18] , \mem[24][17] ,
         \mem[24][16] , \mem[24][15] , \mem[24][14] , \mem[24][13] ,
         \mem[24][12] , \mem[24][11] , \mem[24][10] , \mem[24][9] ,
         \mem[24][8] , \mem[24][7] , \mem[24][6] , \mem[24][5] , \mem[24][4] ,
         \mem[24][3] , \mem[24][2] , \mem[24][1] , \mem[24][0] , \mem[25][23] ,
         \mem[25][22] , \mem[25][21] , \mem[25][20] , \mem[25][19] ,
         \mem[25][18] , \mem[25][17] , \mem[25][16] , \mem[25][15] ,
         \mem[25][14] , \mem[25][13] , \mem[25][12] , \mem[25][11] ,
         \mem[25][10] , \mem[25][9] , \mem[25][8] , \mem[25][7] , \mem[25][6] ,
         \mem[25][5] , \mem[25][4] , \mem[25][3] , \mem[25][2] , \mem[25][1] ,
         \mem[25][0] , \mem[26][23] , \mem[26][22] , \mem[26][21] ,
         \mem[26][20] , \mem[26][19] , \mem[26][18] , \mem[26][17] ,
         \mem[26][16] , \mem[26][15] , \mem[26][14] , \mem[26][13] ,
         \mem[26][12] , \mem[26][11] , \mem[26][10] , \mem[26][9] ,
         \mem[26][8] , \mem[26][7] , \mem[26][6] , \mem[26][5] , \mem[26][4] ,
         \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] , \mem[27][23] ,
         \mem[27][22] , \mem[27][21] , \mem[27][20] , \mem[27][19] ,
         \mem[27][18] , \mem[27][17] , \mem[27][16] , \mem[27][15] ,
         \mem[27][14] , \mem[27][13] , \mem[27][12] , \mem[27][11] ,
         \mem[27][10] , \mem[27][9] , \mem[27][8] , \mem[27][7] , \mem[27][6] ,
         \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] , \mem[27][1] ,
         \mem[27][0] , \mem[28][23] , \mem[28][22] , \mem[28][21] ,
         \mem[28][20] , \mem[28][19] , \mem[28][18] , \mem[28][17] ,
         \mem[28][16] , \mem[28][15] , \mem[28][14] , \mem[28][13] ,
         \mem[28][12] , \mem[28][11] , \mem[28][10] , \mem[28][9] ,
         \mem[28][8] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[29][23] ,
         \mem[29][22] , \mem[29][21] , \mem[29][20] , \mem[29][19] ,
         \mem[29][18] , \mem[29][17] , \mem[29][16] , \mem[29][15] ,
         \mem[29][14] , \mem[29][13] , \mem[29][12] , \mem[29][11] ,
         \mem[29][10] , \mem[29][9] , \mem[29][8] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[30][23] , \mem[30][22] , \mem[30][21] ,
         \mem[30][20] , \mem[30][19] , \mem[30][18] , \mem[30][17] ,
         \mem[30][16] , \mem[30][15] , \mem[30][14] , \mem[30][13] ,
         \mem[30][12] , \mem[30][11] , \mem[30][10] , \mem[30][9] ,
         \mem[30][8] , \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] ,
         \mem[30][3] , \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[31][23] ,
         \mem[31][22] , \mem[31][21] , \mem[31][20] , \mem[31][19] ,
         \mem[31][18] , \mem[31][17] , \mem[31][16] , \mem[31][15] ,
         \mem[31][14] , \mem[31][13] , \mem[31][12] , \mem[31][11] ,
         \mem[31][10] , \mem[31][9] , \mem[31][8] , \mem[31][7] , \mem[31][6] ,
         \mem[31][5] , \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] ,
         \mem[31][0] , n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1938, n1939;

  DFQD1 \mem_reg[0][23]  ( .D(n1937), .CP(clk), .Q(\mem[0][23] ) );
  DFQD1 \mem_reg[0][22]  ( .D(n1936), .CP(clk), .Q(\mem[0][22] ) );
  DFQD1 \mem_reg[0][21]  ( .D(n1935), .CP(clk), .Q(\mem[0][21] ) );
  DFQD1 \mem_reg[0][20]  ( .D(n1934), .CP(clk), .Q(\mem[0][20] ) );
  DFQD1 \mem_reg[0][19]  ( .D(n1933), .CP(clk), .Q(\mem[0][19] ) );
  DFQD1 \mem_reg[0][18]  ( .D(n1932), .CP(clk), .Q(\mem[0][18] ) );
  DFQD1 \mem_reg[0][17]  ( .D(n1931), .CP(clk), .Q(\mem[0][17] ) );
  DFQD1 \mem_reg[0][16]  ( .D(n1930), .CP(clk), .Q(\mem[0][16] ) );
  DFQD1 \mem_reg[0][15]  ( .D(n1929), .CP(clk), .Q(\mem[0][15] ) );
  DFQD1 \mem_reg[0][14]  ( .D(n1928), .CP(clk), .Q(\mem[0][14] ) );
  DFQD1 \mem_reg[0][13]  ( .D(n1927), .CP(clk), .Q(\mem[0][13] ) );
  DFQD1 \mem_reg[0][12]  ( .D(n1926), .CP(clk), .Q(\mem[0][12] ) );
  DFQD1 \mem_reg[0][11]  ( .D(n1925), .CP(clk), .Q(\mem[0][11] ) );
  DFQD1 \mem_reg[0][10]  ( .D(n1924), .CP(clk), .Q(\mem[0][10] ) );
  DFQD1 \mem_reg[0][9]  ( .D(n1923), .CP(clk), .Q(\mem[0][9] ) );
  DFQD1 \mem_reg[0][8]  ( .D(n1922), .CP(clk), .Q(\mem[0][8] ) );
  DFQD1 \mem_reg[0][7]  ( .D(n1921), .CP(clk), .Q(\mem[0][7] ) );
  DFQD1 \mem_reg[0][6]  ( .D(n1920), .CP(clk), .Q(\mem[0][6] ) );
  DFQD1 \mem_reg[0][5]  ( .D(n1919), .CP(clk), .Q(\mem[0][5] ) );
  DFQD1 \mem_reg[0][4]  ( .D(n1918), .CP(clk), .Q(\mem[0][4] ) );
  DFQD1 \mem_reg[0][3]  ( .D(n1917), .CP(clk), .Q(\mem[0][3] ) );
  DFQD1 \mem_reg[0][2]  ( .D(n1916), .CP(clk), .Q(\mem[0][2] ) );
  DFQD1 \mem_reg[0][1]  ( .D(n1915), .CP(clk), .Q(\mem[0][1] ) );
  DFQD1 \mem_reg[0][0]  ( .D(n1914), .CP(clk), .Q(\mem[0][0] ) );
  DFQD1 \mem_reg[1][23]  ( .D(n1913), .CP(clk), .Q(\mem[1][23] ) );
  DFQD1 \mem_reg[1][22]  ( .D(n1912), .CP(clk), .Q(\mem[1][22] ) );
  DFQD1 \mem_reg[1][21]  ( .D(n1911), .CP(clk), .Q(\mem[1][21] ) );
  DFQD1 \mem_reg[1][20]  ( .D(n1910), .CP(clk), .Q(\mem[1][20] ) );
  DFQD1 \mem_reg[1][19]  ( .D(n1909), .CP(clk), .Q(\mem[1][19] ) );
  DFQD1 \mem_reg[1][18]  ( .D(n1908), .CP(clk), .Q(\mem[1][18] ) );
  DFQD1 \mem_reg[1][17]  ( .D(n1907), .CP(clk), .Q(\mem[1][17] ) );
  DFQD1 \mem_reg[1][16]  ( .D(n1906), .CP(clk), .Q(\mem[1][16] ) );
  DFQD1 \mem_reg[1][15]  ( .D(n1905), .CP(clk), .Q(\mem[1][15] ) );
  DFQD1 \mem_reg[1][14]  ( .D(n1904), .CP(clk), .Q(\mem[1][14] ) );
  DFQD1 \mem_reg[1][13]  ( .D(n1903), .CP(clk), .Q(\mem[1][13] ) );
  DFQD1 \mem_reg[1][12]  ( .D(n1902), .CP(clk), .Q(\mem[1][12] ) );
  DFQD1 \mem_reg[1][11]  ( .D(n1901), .CP(clk), .Q(\mem[1][11] ) );
  DFQD1 \mem_reg[1][10]  ( .D(n1900), .CP(clk), .Q(\mem[1][10] ) );
  DFQD1 \mem_reg[1][9]  ( .D(n1899), .CP(clk), .Q(\mem[1][9] ) );
  DFQD1 \mem_reg[1][8]  ( .D(n1898), .CP(clk), .Q(\mem[1][8] ) );
  DFQD1 \mem_reg[1][7]  ( .D(n1897), .CP(clk), .Q(\mem[1][7] ) );
  DFQD1 \mem_reg[1][6]  ( .D(n1896), .CP(clk), .Q(\mem[1][6] ) );
  DFQD1 \mem_reg[1][5]  ( .D(n1895), .CP(clk), .Q(\mem[1][5] ) );
  DFQD1 \mem_reg[1][4]  ( .D(n1894), .CP(clk), .Q(\mem[1][4] ) );
  DFQD1 \mem_reg[1][3]  ( .D(n1893), .CP(clk), .Q(\mem[1][3] ) );
  DFQD1 \mem_reg[1][2]  ( .D(n1892), .CP(clk), .Q(\mem[1][2] ) );
  DFQD1 \mem_reg[1][1]  ( .D(n1891), .CP(clk), .Q(\mem[1][1] ) );
  DFQD1 \mem_reg[1][0]  ( .D(n1890), .CP(clk), .Q(\mem[1][0] ) );
  DFQD1 \mem_reg[2][23]  ( .D(n1889), .CP(clk), .Q(\mem[2][23] ) );
  DFQD1 \mem_reg[2][22]  ( .D(n1888), .CP(clk), .Q(\mem[2][22] ) );
  DFQD1 \mem_reg[2][21]  ( .D(n1887), .CP(clk), .Q(\mem[2][21] ) );
  DFQD1 \mem_reg[2][20]  ( .D(n1886), .CP(clk), .Q(\mem[2][20] ) );
  DFQD1 \mem_reg[2][19]  ( .D(n1885), .CP(clk), .Q(\mem[2][19] ) );
  DFQD1 \mem_reg[2][18]  ( .D(n1884), .CP(clk), .Q(\mem[2][18] ) );
  DFQD1 \mem_reg[2][17]  ( .D(n1883), .CP(clk), .Q(\mem[2][17] ) );
  DFQD1 \mem_reg[2][16]  ( .D(n1882), .CP(clk), .Q(\mem[2][16] ) );
  DFQD1 \mem_reg[2][15]  ( .D(n1881), .CP(clk), .Q(\mem[2][15] ) );
  DFQD1 \mem_reg[2][14]  ( .D(n1880), .CP(clk), .Q(\mem[2][14] ) );
  DFQD1 \mem_reg[2][13]  ( .D(n1879), .CP(clk), .Q(\mem[2][13] ) );
  DFQD1 \mem_reg[2][12]  ( .D(n1878), .CP(clk), .Q(\mem[2][12] ) );
  DFQD1 \mem_reg[2][11]  ( .D(n1877), .CP(clk), .Q(\mem[2][11] ) );
  DFQD1 \mem_reg[2][10]  ( .D(n1876), .CP(clk), .Q(\mem[2][10] ) );
  DFQD1 \mem_reg[2][9]  ( .D(n1875), .CP(clk), .Q(\mem[2][9] ) );
  DFQD1 \mem_reg[2][8]  ( .D(n1874), .CP(clk), .Q(\mem[2][8] ) );
  DFQD1 \mem_reg[2][7]  ( .D(n1873), .CP(clk), .Q(\mem[2][7] ) );
  DFQD1 \mem_reg[2][6]  ( .D(n1872), .CP(clk), .Q(\mem[2][6] ) );
  DFQD1 \mem_reg[2][5]  ( .D(n1871), .CP(clk), .Q(\mem[2][5] ) );
  DFQD1 \mem_reg[2][4]  ( .D(n1870), .CP(clk), .Q(\mem[2][4] ) );
  DFQD1 \mem_reg[2][3]  ( .D(n1869), .CP(clk), .Q(\mem[2][3] ) );
  DFQD1 \mem_reg[2][2]  ( .D(n1868), .CP(clk), .Q(\mem[2][2] ) );
  DFQD1 \mem_reg[2][1]  ( .D(n1867), .CP(clk), .Q(\mem[2][1] ) );
  DFQD1 \mem_reg[2][0]  ( .D(n1866), .CP(clk), .Q(\mem[2][0] ) );
  DFQD1 \mem_reg[3][23]  ( .D(n1865), .CP(clk), .Q(\mem[3][23] ) );
  DFQD1 \mem_reg[3][22]  ( .D(n1864), .CP(clk), .Q(\mem[3][22] ) );
  DFQD1 \mem_reg[3][21]  ( .D(n1863), .CP(clk), .Q(\mem[3][21] ) );
  DFQD1 \mem_reg[3][20]  ( .D(n1862), .CP(clk), .Q(\mem[3][20] ) );
  DFQD1 \mem_reg[3][19]  ( .D(n1861), .CP(clk), .Q(\mem[3][19] ) );
  DFQD1 \mem_reg[3][18]  ( .D(n1860), .CP(clk), .Q(\mem[3][18] ) );
  DFQD1 \mem_reg[3][17]  ( .D(n1859), .CP(clk), .Q(\mem[3][17] ) );
  DFQD1 \mem_reg[3][16]  ( .D(n1858), .CP(clk), .Q(\mem[3][16] ) );
  DFQD1 \mem_reg[3][15]  ( .D(n1857), .CP(clk), .Q(\mem[3][15] ) );
  DFQD1 \mem_reg[3][14]  ( .D(n1856), .CP(clk), .Q(\mem[3][14] ) );
  DFQD1 \mem_reg[3][13]  ( .D(n1855), .CP(clk), .Q(\mem[3][13] ) );
  DFQD1 \mem_reg[3][12]  ( .D(n1854), .CP(clk), .Q(\mem[3][12] ) );
  DFQD1 \mem_reg[3][11]  ( .D(n1853), .CP(clk), .Q(\mem[3][11] ) );
  DFQD1 \mem_reg[3][10]  ( .D(n1852), .CP(clk), .Q(\mem[3][10] ) );
  DFQD1 \mem_reg[3][9]  ( .D(n1851), .CP(clk), .Q(\mem[3][9] ) );
  DFQD1 \mem_reg[3][8]  ( .D(n1850), .CP(clk), .Q(\mem[3][8] ) );
  DFQD1 \mem_reg[3][7]  ( .D(n1849), .CP(clk), .Q(\mem[3][7] ) );
  DFQD1 \mem_reg[3][6]  ( .D(n1848), .CP(clk), .Q(\mem[3][6] ) );
  DFQD1 \mem_reg[3][5]  ( .D(n1847), .CP(clk), .Q(\mem[3][5] ) );
  DFQD1 \mem_reg[3][4]  ( .D(n1846), .CP(clk), .Q(\mem[3][4] ) );
  DFQD1 \mem_reg[3][3]  ( .D(n1845), .CP(clk), .Q(\mem[3][3] ) );
  DFQD1 \mem_reg[3][2]  ( .D(n1844), .CP(clk), .Q(\mem[3][2] ) );
  DFQD1 \mem_reg[3][1]  ( .D(n1843), .CP(clk), .Q(\mem[3][1] ) );
  DFQD1 \mem_reg[3][0]  ( .D(n1842), .CP(clk), .Q(\mem[3][0] ) );
  DFQD1 \mem_reg[4][23]  ( .D(n1841), .CP(clk), .Q(\mem[4][23] ) );
  DFQD1 \mem_reg[4][22]  ( .D(n1840), .CP(clk), .Q(\mem[4][22] ) );
  DFQD1 \mem_reg[4][21]  ( .D(n1839), .CP(clk), .Q(\mem[4][21] ) );
  DFQD1 \mem_reg[4][20]  ( .D(n1838), .CP(clk), .Q(\mem[4][20] ) );
  DFQD1 \mem_reg[4][19]  ( .D(n1837), .CP(clk), .Q(\mem[4][19] ) );
  DFQD1 \mem_reg[4][18]  ( .D(n1836), .CP(clk), .Q(\mem[4][18] ) );
  DFQD1 \mem_reg[4][17]  ( .D(n1835), .CP(clk), .Q(\mem[4][17] ) );
  DFQD1 \mem_reg[4][16]  ( .D(n1834), .CP(clk), .Q(\mem[4][16] ) );
  DFQD1 \mem_reg[4][15]  ( .D(n1833), .CP(clk), .Q(\mem[4][15] ) );
  DFQD1 \mem_reg[4][14]  ( .D(n1832), .CP(clk), .Q(\mem[4][14] ) );
  DFQD1 \mem_reg[4][13]  ( .D(n1831), .CP(clk), .Q(\mem[4][13] ) );
  DFQD1 \mem_reg[4][12]  ( .D(n1830), .CP(clk), .Q(\mem[4][12] ) );
  DFQD1 \mem_reg[4][11]  ( .D(n1829), .CP(clk), .Q(\mem[4][11] ) );
  DFQD1 \mem_reg[4][10]  ( .D(n1828), .CP(clk), .Q(\mem[4][10] ) );
  DFQD1 \mem_reg[4][9]  ( .D(n1827), .CP(clk), .Q(\mem[4][9] ) );
  DFQD1 \mem_reg[4][8]  ( .D(n1826), .CP(clk), .Q(\mem[4][8] ) );
  DFQD1 \mem_reg[4][7]  ( .D(n1825), .CP(clk), .Q(\mem[4][7] ) );
  DFQD1 \mem_reg[4][6]  ( .D(n1824), .CP(clk), .Q(\mem[4][6] ) );
  DFQD1 \mem_reg[4][5]  ( .D(n1823), .CP(clk), .Q(\mem[4][5] ) );
  DFQD1 \mem_reg[4][4]  ( .D(n1822), .CP(clk), .Q(\mem[4][4] ) );
  DFQD1 \mem_reg[4][3]  ( .D(n1821), .CP(clk), .Q(\mem[4][3] ) );
  DFQD1 \mem_reg[4][2]  ( .D(n1820), .CP(clk), .Q(\mem[4][2] ) );
  DFQD1 \mem_reg[4][1]  ( .D(n1819), .CP(clk), .Q(\mem[4][1] ) );
  DFQD1 \mem_reg[4][0]  ( .D(n1818), .CP(clk), .Q(\mem[4][0] ) );
  DFQD1 \mem_reg[5][23]  ( .D(n1817), .CP(clk), .Q(\mem[5][23] ) );
  DFQD1 \mem_reg[5][22]  ( .D(n1816), .CP(clk), .Q(\mem[5][22] ) );
  DFQD1 \mem_reg[5][21]  ( .D(n1815), .CP(clk), .Q(\mem[5][21] ) );
  DFQD1 \mem_reg[5][20]  ( .D(n1814), .CP(clk), .Q(\mem[5][20] ) );
  DFQD1 \mem_reg[5][19]  ( .D(n1813), .CP(clk), .Q(\mem[5][19] ) );
  DFQD1 \mem_reg[5][18]  ( .D(n1812), .CP(clk), .Q(\mem[5][18] ) );
  DFQD1 \mem_reg[5][17]  ( .D(n1811), .CP(clk), .Q(\mem[5][17] ) );
  DFQD1 \mem_reg[5][16]  ( .D(n1810), .CP(clk), .Q(\mem[5][16] ) );
  DFQD1 \mem_reg[5][15]  ( .D(n1809), .CP(clk), .Q(\mem[5][15] ) );
  DFQD1 \mem_reg[5][14]  ( .D(n1808), .CP(clk), .Q(\mem[5][14] ) );
  DFQD1 \mem_reg[5][13]  ( .D(n1807), .CP(clk), .Q(\mem[5][13] ) );
  DFQD1 \mem_reg[5][12]  ( .D(n1806), .CP(clk), .Q(\mem[5][12] ) );
  DFQD1 \mem_reg[5][11]  ( .D(n1805), .CP(clk), .Q(\mem[5][11] ) );
  DFQD1 \mem_reg[5][10]  ( .D(n1804), .CP(clk), .Q(\mem[5][10] ) );
  DFQD1 \mem_reg[5][9]  ( .D(n1803), .CP(clk), .Q(\mem[5][9] ) );
  DFQD1 \mem_reg[5][8]  ( .D(n1802), .CP(clk), .Q(\mem[5][8] ) );
  DFQD1 \mem_reg[5][7]  ( .D(n1801), .CP(clk), .Q(\mem[5][7] ) );
  DFQD1 \mem_reg[5][6]  ( .D(n1800), .CP(clk), .Q(\mem[5][6] ) );
  DFQD1 \mem_reg[5][5]  ( .D(n1799), .CP(clk), .Q(\mem[5][5] ) );
  DFQD1 \mem_reg[5][4]  ( .D(n1798), .CP(clk), .Q(\mem[5][4] ) );
  DFQD1 \mem_reg[5][3]  ( .D(n1797), .CP(clk), .Q(\mem[5][3] ) );
  DFQD1 \mem_reg[5][2]  ( .D(n1796), .CP(clk), .Q(\mem[5][2] ) );
  DFQD1 \mem_reg[5][1]  ( .D(n1795), .CP(clk), .Q(\mem[5][1] ) );
  DFQD1 \mem_reg[5][0]  ( .D(n1794), .CP(clk), .Q(\mem[5][0] ) );
  DFQD1 \mem_reg[6][23]  ( .D(n1793), .CP(clk), .Q(\mem[6][23] ) );
  DFQD1 \mem_reg[6][22]  ( .D(n1792), .CP(clk), .Q(\mem[6][22] ) );
  DFQD1 \mem_reg[6][21]  ( .D(n1791), .CP(clk), .Q(\mem[6][21] ) );
  DFQD1 \mem_reg[6][20]  ( .D(n1790), .CP(clk), .Q(\mem[6][20] ) );
  DFQD1 \mem_reg[6][19]  ( .D(n1789), .CP(clk), .Q(\mem[6][19] ) );
  DFQD1 \mem_reg[6][18]  ( .D(n1788), .CP(clk), .Q(\mem[6][18] ) );
  DFQD1 \mem_reg[6][17]  ( .D(n1787), .CP(clk), .Q(\mem[6][17] ) );
  DFQD1 \mem_reg[6][16]  ( .D(n1786), .CP(clk), .Q(\mem[6][16] ) );
  DFQD1 \mem_reg[6][15]  ( .D(n1785), .CP(clk), .Q(\mem[6][15] ) );
  DFQD1 \mem_reg[6][14]  ( .D(n1784), .CP(clk), .Q(\mem[6][14] ) );
  DFQD1 \mem_reg[6][13]  ( .D(n1783), .CP(clk), .Q(\mem[6][13] ) );
  DFQD1 \mem_reg[6][12]  ( .D(n1782), .CP(clk), .Q(\mem[6][12] ) );
  DFQD1 \mem_reg[6][11]  ( .D(n1781), .CP(clk), .Q(\mem[6][11] ) );
  DFQD1 \mem_reg[6][10]  ( .D(n1780), .CP(clk), .Q(\mem[6][10] ) );
  DFQD1 \mem_reg[6][9]  ( .D(n1779), .CP(clk), .Q(\mem[6][9] ) );
  DFQD1 \mem_reg[6][8]  ( .D(n1778), .CP(clk), .Q(\mem[6][8] ) );
  DFQD1 \mem_reg[6][7]  ( .D(n1777), .CP(clk), .Q(\mem[6][7] ) );
  DFQD1 \mem_reg[6][6]  ( .D(n1776), .CP(clk), .Q(\mem[6][6] ) );
  DFQD1 \mem_reg[6][5]  ( .D(n1775), .CP(clk), .Q(\mem[6][5] ) );
  DFQD1 \mem_reg[6][4]  ( .D(n1774), .CP(clk), .Q(\mem[6][4] ) );
  DFQD1 \mem_reg[6][3]  ( .D(n1773), .CP(clk), .Q(\mem[6][3] ) );
  DFQD1 \mem_reg[6][2]  ( .D(n1772), .CP(clk), .Q(\mem[6][2] ) );
  DFQD1 \mem_reg[6][1]  ( .D(n1771), .CP(clk), .Q(\mem[6][1] ) );
  DFQD1 \mem_reg[6][0]  ( .D(n1770), .CP(clk), .Q(\mem[6][0] ) );
  DFQD1 \mem_reg[7][23]  ( .D(n1769), .CP(clk), .Q(\mem[7][23] ) );
  DFQD1 \mem_reg[7][22]  ( .D(n1768), .CP(clk), .Q(\mem[7][22] ) );
  DFQD1 \mem_reg[7][21]  ( .D(n1767), .CP(clk), .Q(\mem[7][21] ) );
  DFQD1 \mem_reg[7][20]  ( .D(n1766), .CP(clk), .Q(\mem[7][20] ) );
  DFQD1 \mem_reg[7][19]  ( .D(n1765), .CP(clk), .Q(\mem[7][19] ) );
  DFQD1 \mem_reg[7][18]  ( .D(n1764), .CP(clk), .Q(\mem[7][18] ) );
  DFQD1 \mem_reg[7][17]  ( .D(n1763), .CP(clk), .Q(\mem[7][17] ) );
  DFQD1 \mem_reg[7][16]  ( .D(n1762), .CP(clk), .Q(\mem[7][16] ) );
  DFQD1 \mem_reg[7][15]  ( .D(n1761), .CP(clk), .Q(\mem[7][15] ) );
  DFQD1 \mem_reg[7][14]  ( .D(n1760), .CP(clk), .Q(\mem[7][14] ) );
  DFQD1 \mem_reg[7][13]  ( .D(n1759), .CP(clk), .Q(\mem[7][13] ) );
  DFQD1 \mem_reg[7][12]  ( .D(n1758), .CP(clk), .Q(\mem[7][12] ) );
  DFQD1 \mem_reg[7][11]  ( .D(n1757), .CP(clk), .Q(\mem[7][11] ) );
  DFQD1 \mem_reg[7][10]  ( .D(n1756), .CP(clk), .Q(\mem[7][10] ) );
  DFQD1 \mem_reg[7][9]  ( .D(n1755), .CP(clk), .Q(\mem[7][9] ) );
  DFQD1 \mem_reg[7][8]  ( .D(n1754), .CP(clk), .Q(\mem[7][8] ) );
  DFQD1 \mem_reg[7][7]  ( .D(n1753), .CP(clk), .Q(\mem[7][7] ) );
  DFQD1 \mem_reg[7][6]  ( .D(n1752), .CP(clk), .Q(\mem[7][6] ) );
  DFQD1 \mem_reg[7][5]  ( .D(n1751), .CP(clk), .Q(\mem[7][5] ) );
  DFQD1 \mem_reg[7][4]  ( .D(n1750), .CP(clk), .Q(\mem[7][4] ) );
  DFQD1 \mem_reg[7][3]  ( .D(n1749), .CP(clk), .Q(\mem[7][3] ) );
  DFQD1 \mem_reg[7][2]  ( .D(n1748), .CP(clk), .Q(\mem[7][2] ) );
  DFQD1 \mem_reg[7][1]  ( .D(n1747), .CP(clk), .Q(\mem[7][1] ) );
  DFQD1 \mem_reg[7][0]  ( .D(n1746), .CP(clk), .Q(\mem[7][0] ) );
  DFQD1 \mem_reg[8][23]  ( .D(n1745), .CP(clk), .Q(\mem[8][23] ) );
  DFQD1 \mem_reg[8][22]  ( .D(n1744), .CP(clk), .Q(\mem[8][22] ) );
  DFQD1 \mem_reg[8][21]  ( .D(n1743), .CP(clk), .Q(\mem[8][21] ) );
  DFQD1 \mem_reg[8][20]  ( .D(n1742), .CP(clk), .Q(\mem[8][20] ) );
  DFQD1 \mem_reg[8][19]  ( .D(n1741), .CP(clk), .Q(\mem[8][19] ) );
  DFQD1 \mem_reg[8][18]  ( .D(n1740), .CP(clk), .Q(\mem[8][18] ) );
  DFQD1 \mem_reg[8][17]  ( .D(n1739), .CP(clk), .Q(\mem[8][17] ) );
  DFQD1 \mem_reg[8][16]  ( .D(n1738), .CP(clk), .Q(\mem[8][16] ) );
  DFQD1 \mem_reg[8][15]  ( .D(n1737), .CP(clk), .Q(\mem[8][15] ) );
  DFQD1 \mem_reg[8][14]  ( .D(n1736), .CP(clk), .Q(\mem[8][14] ) );
  DFQD1 \mem_reg[8][13]  ( .D(n1735), .CP(clk), .Q(\mem[8][13] ) );
  DFQD1 \mem_reg[8][12]  ( .D(n1734), .CP(clk), .Q(\mem[8][12] ) );
  DFQD1 \mem_reg[8][11]  ( .D(n1733), .CP(clk), .Q(\mem[8][11] ) );
  DFQD1 \mem_reg[8][10]  ( .D(n1732), .CP(clk), .Q(\mem[8][10] ) );
  DFQD1 \mem_reg[8][9]  ( .D(n1731), .CP(clk), .Q(\mem[8][9] ) );
  DFQD1 \mem_reg[8][8]  ( .D(n1730), .CP(clk), .Q(\mem[8][8] ) );
  DFQD1 \mem_reg[8][7]  ( .D(n1729), .CP(clk), .Q(\mem[8][7] ) );
  DFQD1 \mem_reg[8][6]  ( .D(n1728), .CP(clk), .Q(\mem[8][6] ) );
  DFQD1 \mem_reg[8][5]  ( .D(n1727), .CP(clk), .Q(\mem[8][5] ) );
  DFQD1 \mem_reg[8][4]  ( .D(n1726), .CP(clk), .Q(\mem[8][4] ) );
  DFQD1 \mem_reg[8][3]  ( .D(n1725), .CP(clk), .Q(\mem[8][3] ) );
  DFQD1 \mem_reg[8][2]  ( .D(n1724), .CP(clk), .Q(\mem[8][2] ) );
  DFQD1 \mem_reg[8][1]  ( .D(n1723), .CP(clk), .Q(\mem[8][1] ) );
  DFQD1 \mem_reg[8][0]  ( .D(n1722), .CP(clk), .Q(\mem[8][0] ) );
  DFQD1 \mem_reg[9][23]  ( .D(n1721), .CP(clk), .Q(\mem[9][23] ) );
  DFQD1 \mem_reg[9][22]  ( .D(n1720), .CP(clk), .Q(\mem[9][22] ) );
  DFQD1 \mem_reg[9][21]  ( .D(n1719), .CP(clk), .Q(\mem[9][21] ) );
  DFQD1 \mem_reg[9][20]  ( .D(n1718), .CP(clk), .Q(\mem[9][20] ) );
  DFQD1 \mem_reg[9][19]  ( .D(n1717), .CP(clk), .Q(\mem[9][19] ) );
  DFQD1 \mem_reg[9][18]  ( .D(n1716), .CP(clk), .Q(\mem[9][18] ) );
  DFQD1 \mem_reg[9][17]  ( .D(n1715), .CP(clk), .Q(\mem[9][17] ) );
  DFQD1 \mem_reg[9][16]  ( .D(n1714), .CP(clk), .Q(\mem[9][16] ) );
  DFQD1 \mem_reg[9][15]  ( .D(n1713), .CP(clk), .Q(\mem[9][15] ) );
  DFQD1 \mem_reg[9][14]  ( .D(n1712), .CP(clk), .Q(\mem[9][14] ) );
  DFQD1 \mem_reg[9][13]  ( .D(n1711), .CP(clk), .Q(\mem[9][13] ) );
  DFQD1 \mem_reg[9][12]  ( .D(n1710), .CP(clk), .Q(\mem[9][12] ) );
  DFQD1 \mem_reg[9][11]  ( .D(n1709), .CP(clk), .Q(\mem[9][11] ) );
  DFQD1 \mem_reg[9][10]  ( .D(n1708), .CP(clk), .Q(\mem[9][10] ) );
  DFQD1 \mem_reg[9][9]  ( .D(n1707), .CP(clk), .Q(\mem[9][9] ) );
  DFQD1 \mem_reg[9][8]  ( .D(n1706), .CP(clk), .Q(\mem[9][8] ) );
  DFQD1 \mem_reg[9][7]  ( .D(n1705), .CP(clk), .Q(\mem[9][7] ) );
  DFQD1 \mem_reg[9][6]  ( .D(n1704), .CP(clk), .Q(\mem[9][6] ) );
  DFQD1 \mem_reg[9][5]  ( .D(n1703), .CP(clk), .Q(\mem[9][5] ) );
  DFQD1 \mem_reg[9][4]  ( .D(n1702), .CP(clk), .Q(\mem[9][4] ) );
  DFQD1 \mem_reg[9][3]  ( .D(n1701), .CP(clk), .Q(\mem[9][3] ) );
  DFQD1 \mem_reg[9][2]  ( .D(n1700), .CP(clk), .Q(\mem[9][2] ) );
  DFQD1 \mem_reg[9][1]  ( .D(n1699), .CP(clk), .Q(\mem[9][1] ) );
  DFQD1 \mem_reg[9][0]  ( .D(n1698), .CP(clk), .Q(\mem[9][0] ) );
  DFQD1 \mem_reg[10][23]  ( .D(n1697), .CP(clk), .Q(\mem[10][23] ) );
  DFQD1 \mem_reg[10][22]  ( .D(n1696), .CP(clk), .Q(\mem[10][22] ) );
  DFQD1 \mem_reg[10][21]  ( .D(n1695), .CP(clk), .Q(\mem[10][21] ) );
  DFQD1 \mem_reg[10][20]  ( .D(n1694), .CP(clk), .Q(\mem[10][20] ) );
  DFQD1 \mem_reg[10][19]  ( .D(n1693), .CP(clk), .Q(\mem[10][19] ) );
  DFQD1 \mem_reg[10][18]  ( .D(n1692), .CP(clk), .Q(\mem[10][18] ) );
  DFQD1 \mem_reg[10][17]  ( .D(n1691), .CP(clk), .Q(\mem[10][17] ) );
  DFQD1 \mem_reg[10][16]  ( .D(n1690), .CP(clk), .Q(\mem[10][16] ) );
  DFQD1 \mem_reg[10][15]  ( .D(n1689), .CP(clk), .Q(\mem[10][15] ) );
  DFQD1 \mem_reg[10][14]  ( .D(n1688), .CP(clk), .Q(\mem[10][14] ) );
  DFQD1 \mem_reg[10][13]  ( .D(n1687), .CP(clk), .Q(\mem[10][13] ) );
  DFQD1 \mem_reg[10][12]  ( .D(n1686), .CP(clk), .Q(\mem[10][12] ) );
  DFQD1 \mem_reg[10][11]  ( .D(n1685), .CP(clk), .Q(\mem[10][11] ) );
  DFQD1 \mem_reg[10][10]  ( .D(n1684), .CP(clk), .Q(\mem[10][10] ) );
  DFQD1 \mem_reg[10][9]  ( .D(n1683), .CP(clk), .Q(\mem[10][9] ) );
  DFQD1 \mem_reg[10][8]  ( .D(n1682), .CP(clk), .Q(\mem[10][8] ) );
  DFQD1 \mem_reg[10][7]  ( .D(n1681), .CP(clk), .Q(\mem[10][7] ) );
  DFQD1 \mem_reg[10][6]  ( .D(n1680), .CP(clk), .Q(\mem[10][6] ) );
  DFQD1 \mem_reg[10][5]  ( .D(n1679), .CP(clk), .Q(\mem[10][5] ) );
  DFQD1 \mem_reg[10][4]  ( .D(n1678), .CP(clk), .Q(\mem[10][4] ) );
  DFQD1 \mem_reg[10][3]  ( .D(n1677), .CP(clk), .Q(\mem[10][3] ) );
  DFQD1 \mem_reg[10][2]  ( .D(n1676), .CP(clk), .Q(\mem[10][2] ) );
  DFQD1 \mem_reg[10][1]  ( .D(n1675), .CP(clk), .Q(\mem[10][1] ) );
  DFQD1 \mem_reg[10][0]  ( .D(n1674), .CP(clk), .Q(\mem[10][0] ) );
  DFQD1 \mem_reg[11][23]  ( .D(n1673), .CP(clk), .Q(\mem[11][23] ) );
  DFQD1 \mem_reg[11][22]  ( .D(n1672), .CP(clk), .Q(\mem[11][22] ) );
  DFQD1 \mem_reg[11][21]  ( .D(n1671), .CP(clk), .Q(\mem[11][21] ) );
  DFQD1 \mem_reg[11][20]  ( .D(n1670), .CP(clk), .Q(\mem[11][20] ) );
  DFQD1 \mem_reg[11][19]  ( .D(n1669), .CP(clk), .Q(\mem[11][19] ) );
  DFQD1 \mem_reg[11][18]  ( .D(n1668), .CP(clk), .Q(\mem[11][18] ) );
  DFQD1 \mem_reg[11][17]  ( .D(n1667), .CP(clk), .Q(\mem[11][17] ) );
  DFQD1 \mem_reg[11][16]  ( .D(n1666), .CP(clk), .Q(\mem[11][16] ) );
  DFQD1 \mem_reg[11][15]  ( .D(n1665), .CP(clk), .Q(\mem[11][15] ) );
  DFQD1 \mem_reg[11][14]  ( .D(n1664), .CP(clk), .Q(\mem[11][14] ) );
  DFQD1 \mem_reg[11][13]  ( .D(n1663), .CP(clk), .Q(\mem[11][13] ) );
  DFQD1 \mem_reg[11][12]  ( .D(n1662), .CP(clk), .Q(\mem[11][12] ) );
  DFQD1 \mem_reg[11][11]  ( .D(n1661), .CP(clk), .Q(\mem[11][11] ) );
  DFQD1 \mem_reg[11][10]  ( .D(n1660), .CP(clk), .Q(\mem[11][10] ) );
  DFQD1 \mem_reg[11][9]  ( .D(n1659), .CP(clk), .Q(\mem[11][9] ) );
  DFQD1 \mem_reg[11][8]  ( .D(n1658), .CP(clk), .Q(\mem[11][8] ) );
  DFQD1 \mem_reg[11][7]  ( .D(n1657), .CP(clk), .Q(\mem[11][7] ) );
  DFQD1 \mem_reg[11][6]  ( .D(n1656), .CP(clk), .Q(\mem[11][6] ) );
  DFQD1 \mem_reg[11][5]  ( .D(n1655), .CP(clk), .Q(\mem[11][5] ) );
  DFQD1 \mem_reg[11][4]  ( .D(n1654), .CP(clk), .Q(\mem[11][4] ) );
  DFQD1 \mem_reg[11][3]  ( .D(n1653), .CP(clk), .Q(\mem[11][3] ) );
  DFQD1 \mem_reg[11][2]  ( .D(n1652), .CP(clk), .Q(\mem[11][2] ) );
  DFQD1 \mem_reg[11][1]  ( .D(n1651), .CP(clk), .Q(\mem[11][1] ) );
  DFQD1 \mem_reg[11][0]  ( .D(n1650), .CP(clk), .Q(\mem[11][0] ) );
  DFQD1 \mem_reg[12][23]  ( .D(n1649), .CP(clk), .Q(\mem[12][23] ) );
  DFQD1 \mem_reg[12][22]  ( .D(n1648), .CP(clk), .Q(\mem[12][22] ) );
  DFQD1 \mem_reg[12][21]  ( .D(n1647), .CP(clk), .Q(\mem[12][21] ) );
  DFQD1 \mem_reg[12][20]  ( .D(n1646), .CP(clk), .Q(\mem[12][20] ) );
  DFQD1 \mem_reg[12][19]  ( .D(n1645), .CP(clk), .Q(\mem[12][19] ) );
  DFQD1 \mem_reg[12][18]  ( .D(n1644), .CP(clk), .Q(\mem[12][18] ) );
  DFQD1 \mem_reg[12][17]  ( .D(n1643), .CP(clk), .Q(\mem[12][17] ) );
  DFQD1 \mem_reg[12][16]  ( .D(n1642), .CP(clk), .Q(\mem[12][16] ) );
  DFQD1 \mem_reg[12][15]  ( .D(n1641), .CP(clk), .Q(\mem[12][15] ) );
  DFQD1 \mem_reg[12][14]  ( .D(n1640), .CP(clk), .Q(\mem[12][14] ) );
  DFQD1 \mem_reg[12][13]  ( .D(n1639), .CP(clk), .Q(\mem[12][13] ) );
  DFQD1 \mem_reg[12][12]  ( .D(n1638), .CP(clk), .Q(\mem[12][12] ) );
  DFQD1 \mem_reg[12][11]  ( .D(n1637), .CP(clk), .Q(\mem[12][11] ) );
  DFQD1 \mem_reg[12][10]  ( .D(n1636), .CP(clk), .Q(\mem[12][10] ) );
  DFQD1 \mem_reg[12][9]  ( .D(n1635), .CP(clk), .Q(\mem[12][9] ) );
  DFQD1 \mem_reg[12][8]  ( .D(n1634), .CP(clk), .Q(\mem[12][8] ) );
  DFQD1 \mem_reg[12][7]  ( .D(n1633), .CP(clk), .Q(\mem[12][7] ) );
  DFQD1 \mem_reg[12][6]  ( .D(n1632), .CP(clk), .Q(\mem[12][6] ) );
  DFQD1 \mem_reg[12][5]  ( .D(n1631), .CP(clk), .Q(\mem[12][5] ) );
  DFQD1 \mem_reg[12][4]  ( .D(n1630), .CP(clk), .Q(\mem[12][4] ) );
  DFQD1 \mem_reg[12][3]  ( .D(n1629), .CP(clk), .Q(\mem[12][3] ) );
  DFQD1 \mem_reg[12][2]  ( .D(n1628), .CP(clk), .Q(\mem[12][2] ) );
  DFQD1 \mem_reg[12][1]  ( .D(n1627), .CP(clk), .Q(\mem[12][1] ) );
  DFQD1 \mem_reg[12][0]  ( .D(n1626), .CP(clk), .Q(\mem[12][0] ) );
  DFQD1 \mem_reg[13][23]  ( .D(n1625), .CP(clk), .Q(\mem[13][23] ) );
  DFQD1 \mem_reg[13][22]  ( .D(n1624), .CP(clk), .Q(\mem[13][22] ) );
  DFQD1 \mem_reg[13][21]  ( .D(n1623), .CP(clk), .Q(\mem[13][21] ) );
  DFQD1 \mem_reg[13][20]  ( .D(n1622), .CP(clk), .Q(\mem[13][20] ) );
  DFQD1 \mem_reg[13][19]  ( .D(n1621), .CP(clk), .Q(\mem[13][19] ) );
  DFQD1 \mem_reg[13][18]  ( .D(n1620), .CP(clk), .Q(\mem[13][18] ) );
  DFQD1 \mem_reg[13][17]  ( .D(n1619), .CP(clk), .Q(\mem[13][17] ) );
  DFQD1 \mem_reg[13][16]  ( .D(n1618), .CP(clk), .Q(\mem[13][16] ) );
  DFQD1 \mem_reg[13][15]  ( .D(n1617), .CP(clk), .Q(\mem[13][15] ) );
  DFQD1 \mem_reg[13][14]  ( .D(n1616), .CP(clk), .Q(\mem[13][14] ) );
  DFQD1 \mem_reg[13][13]  ( .D(n1615), .CP(clk), .Q(\mem[13][13] ) );
  DFQD1 \mem_reg[13][12]  ( .D(n1614), .CP(clk), .Q(\mem[13][12] ) );
  DFQD1 \mem_reg[13][11]  ( .D(n1613), .CP(clk), .Q(\mem[13][11] ) );
  DFQD1 \mem_reg[13][10]  ( .D(n1612), .CP(clk), .Q(\mem[13][10] ) );
  DFQD1 \mem_reg[13][9]  ( .D(n1611), .CP(clk), .Q(\mem[13][9] ) );
  DFQD1 \mem_reg[13][8]  ( .D(n1610), .CP(clk), .Q(\mem[13][8] ) );
  DFQD1 \mem_reg[13][7]  ( .D(n1609), .CP(clk), .Q(\mem[13][7] ) );
  DFQD1 \mem_reg[13][6]  ( .D(n1608), .CP(clk), .Q(\mem[13][6] ) );
  DFQD1 \mem_reg[13][5]  ( .D(n1607), .CP(clk), .Q(\mem[13][5] ) );
  DFQD1 \mem_reg[13][4]  ( .D(n1606), .CP(clk), .Q(\mem[13][4] ) );
  DFQD1 \mem_reg[13][3]  ( .D(n1605), .CP(clk), .Q(\mem[13][3] ) );
  DFQD1 \mem_reg[13][2]  ( .D(n1604), .CP(clk), .Q(\mem[13][2] ) );
  DFQD1 \mem_reg[13][1]  ( .D(n1603), .CP(clk), .Q(\mem[13][1] ) );
  DFQD1 \mem_reg[13][0]  ( .D(n1602), .CP(clk), .Q(\mem[13][0] ) );
  DFQD1 \mem_reg[14][23]  ( .D(n1601), .CP(clk), .Q(\mem[14][23] ) );
  DFQD1 \mem_reg[14][22]  ( .D(n1600), .CP(clk), .Q(\mem[14][22] ) );
  DFQD1 \mem_reg[14][21]  ( .D(n1599), .CP(clk), .Q(\mem[14][21] ) );
  DFQD1 \mem_reg[14][20]  ( .D(n1598), .CP(clk), .Q(\mem[14][20] ) );
  DFQD1 \mem_reg[14][19]  ( .D(n1597), .CP(clk), .Q(\mem[14][19] ) );
  DFQD1 \mem_reg[14][18]  ( .D(n1596), .CP(clk), .Q(\mem[14][18] ) );
  DFQD1 \mem_reg[14][17]  ( .D(n1595), .CP(clk), .Q(\mem[14][17] ) );
  DFQD1 \mem_reg[14][16]  ( .D(n1594), .CP(clk), .Q(\mem[14][16] ) );
  DFQD1 \mem_reg[14][15]  ( .D(n1593), .CP(clk), .Q(\mem[14][15] ) );
  DFQD1 \mem_reg[14][14]  ( .D(n1592), .CP(clk), .Q(\mem[14][14] ) );
  DFQD1 \mem_reg[14][13]  ( .D(n1591), .CP(clk), .Q(\mem[14][13] ) );
  DFQD1 \mem_reg[14][12]  ( .D(n1590), .CP(clk), .Q(\mem[14][12] ) );
  DFQD1 \mem_reg[14][11]  ( .D(n1589), .CP(clk), .Q(\mem[14][11] ) );
  DFQD1 \mem_reg[14][10]  ( .D(n1588), .CP(clk), .Q(\mem[14][10] ) );
  DFQD1 \mem_reg[14][9]  ( .D(n1587), .CP(clk), .Q(\mem[14][9] ) );
  DFQD1 \mem_reg[14][8]  ( .D(n1586), .CP(clk), .Q(\mem[14][8] ) );
  DFQD1 \mem_reg[14][7]  ( .D(n1585), .CP(clk), .Q(\mem[14][7] ) );
  DFQD1 \mem_reg[14][6]  ( .D(n1584), .CP(clk), .Q(\mem[14][6] ) );
  DFQD1 \mem_reg[14][5]  ( .D(n1583), .CP(clk), .Q(\mem[14][5] ) );
  DFQD1 \mem_reg[14][4]  ( .D(n1582), .CP(clk), .Q(\mem[14][4] ) );
  DFQD1 \mem_reg[14][3]  ( .D(n1581), .CP(clk), .Q(\mem[14][3] ) );
  DFQD1 \mem_reg[14][2]  ( .D(n1580), .CP(clk), .Q(\mem[14][2] ) );
  DFQD1 \mem_reg[14][1]  ( .D(n1579), .CP(clk), .Q(\mem[14][1] ) );
  DFQD1 \mem_reg[14][0]  ( .D(n1578), .CP(clk), .Q(\mem[14][0] ) );
  DFQD1 \mem_reg[15][23]  ( .D(n1577), .CP(clk), .Q(\mem[15][23] ) );
  DFQD1 \mem_reg[15][22]  ( .D(n1576), .CP(clk), .Q(\mem[15][22] ) );
  DFQD1 \mem_reg[15][21]  ( .D(n1575), .CP(clk), .Q(\mem[15][21] ) );
  DFQD1 \mem_reg[15][20]  ( .D(n1574), .CP(clk), .Q(\mem[15][20] ) );
  DFQD1 \mem_reg[15][19]  ( .D(n1573), .CP(clk), .Q(\mem[15][19] ) );
  DFQD1 \mem_reg[15][18]  ( .D(n1572), .CP(clk), .Q(\mem[15][18] ) );
  DFQD1 \mem_reg[15][17]  ( .D(n1571), .CP(clk), .Q(\mem[15][17] ) );
  DFQD1 \mem_reg[15][16]  ( .D(n1570), .CP(clk), .Q(\mem[15][16] ) );
  DFQD1 \mem_reg[15][15]  ( .D(n1569), .CP(clk), .Q(\mem[15][15] ) );
  DFQD1 \mem_reg[15][14]  ( .D(n1568), .CP(clk), .Q(\mem[15][14] ) );
  DFQD1 \mem_reg[15][13]  ( .D(n1567), .CP(clk), .Q(\mem[15][13] ) );
  DFQD1 \mem_reg[15][12]  ( .D(n1566), .CP(clk), .Q(\mem[15][12] ) );
  DFQD1 \mem_reg[15][11]  ( .D(n1565), .CP(clk), .Q(\mem[15][11] ) );
  DFQD1 \mem_reg[15][10]  ( .D(n1564), .CP(clk), .Q(\mem[15][10] ) );
  DFQD1 \mem_reg[15][9]  ( .D(n1563), .CP(clk), .Q(\mem[15][9] ) );
  DFQD1 \mem_reg[15][8]  ( .D(n1562), .CP(clk), .Q(\mem[15][8] ) );
  DFQD1 \mem_reg[15][7]  ( .D(n1561), .CP(clk), .Q(\mem[15][7] ) );
  DFQD1 \mem_reg[15][6]  ( .D(n1560), .CP(clk), .Q(\mem[15][6] ) );
  DFQD1 \mem_reg[15][5]  ( .D(n1559), .CP(clk), .Q(\mem[15][5] ) );
  DFQD1 \mem_reg[15][4]  ( .D(n1558), .CP(clk), .Q(\mem[15][4] ) );
  DFQD1 \mem_reg[15][3]  ( .D(n1557), .CP(clk), .Q(\mem[15][3] ) );
  DFQD1 \mem_reg[15][2]  ( .D(n1556), .CP(clk), .Q(\mem[15][2] ) );
  DFQD1 \mem_reg[15][1]  ( .D(n1555), .CP(clk), .Q(\mem[15][1] ) );
  DFQD1 \mem_reg[15][0]  ( .D(n1554), .CP(clk), .Q(\mem[15][0] ) );
  DFQD1 \mem_reg[16][23]  ( .D(n1553), .CP(clk), .Q(\mem[16][23] ) );
  DFQD1 \mem_reg[16][22]  ( .D(n1552), .CP(clk), .Q(\mem[16][22] ) );
  DFQD1 \mem_reg[16][21]  ( .D(n1551), .CP(clk), .Q(\mem[16][21] ) );
  DFQD1 \mem_reg[16][20]  ( .D(n1550), .CP(clk), .Q(\mem[16][20] ) );
  DFQD1 \mem_reg[16][19]  ( .D(n1549), .CP(clk), .Q(\mem[16][19] ) );
  DFQD1 \mem_reg[16][18]  ( .D(n1548), .CP(clk), .Q(\mem[16][18] ) );
  DFQD1 \mem_reg[16][17]  ( .D(n1547), .CP(clk), .Q(\mem[16][17] ) );
  DFQD1 \mem_reg[16][16]  ( .D(n1546), .CP(clk), .Q(\mem[16][16] ) );
  DFQD1 \mem_reg[16][15]  ( .D(n1545), .CP(clk), .Q(\mem[16][15] ) );
  DFQD1 \mem_reg[16][14]  ( .D(n1544), .CP(clk), .Q(\mem[16][14] ) );
  DFQD1 \mem_reg[16][13]  ( .D(n1543), .CP(clk), .Q(\mem[16][13] ) );
  DFQD1 \mem_reg[16][12]  ( .D(n1542), .CP(clk), .Q(\mem[16][12] ) );
  DFQD1 \mem_reg[16][11]  ( .D(n1541), .CP(clk), .Q(\mem[16][11] ) );
  DFQD1 \mem_reg[16][10]  ( .D(n1540), .CP(clk), .Q(\mem[16][10] ) );
  DFQD1 \mem_reg[16][9]  ( .D(n1539), .CP(clk), .Q(\mem[16][9] ) );
  DFQD1 \mem_reg[16][8]  ( .D(n1538), .CP(clk), .Q(\mem[16][8] ) );
  DFQD1 \mem_reg[16][7]  ( .D(n1537), .CP(clk), .Q(\mem[16][7] ) );
  DFQD1 \mem_reg[16][6]  ( .D(n1536), .CP(clk), .Q(\mem[16][6] ) );
  DFQD1 \mem_reg[16][5]  ( .D(n1535), .CP(clk), .Q(\mem[16][5] ) );
  DFQD1 \mem_reg[16][4]  ( .D(n1534), .CP(clk), .Q(\mem[16][4] ) );
  DFQD1 \mem_reg[16][3]  ( .D(n1533), .CP(clk), .Q(\mem[16][3] ) );
  DFQD1 \mem_reg[16][2]  ( .D(n1532), .CP(clk), .Q(\mem[16][2] ) );
  DFQD1 \mem_reg[16][1]  ( .D(n1531), .CP(clk), .Q(\mem[16][1] ) );
  DFQD1 \mem_reg[16][0]  ( .D(n1530), .CP(clk), .Q(\mem[16][0] ) );
  DFQD1 \mem_reg[17][23]  ( .D(n1529), .CP(clk), .Q(\mem[17][23] ) );
  DFQD1 \mem_reg[17][22]  ( .D(n1528), .CP(clk), .Q(\mem[17][22] ) );
  DFQD1 \mem_reg[17][21]  ( .D(n1527), .CP(clk), .Q(\mem[17][21] ) );
  DFQD1 \mem_reg[17][20]  ( .D(n1526), .CP(clk), .Q(\mem[17][20] ) );
  DFQD1 \mem_reg[17][19]  ( .D(n1525), .CP(clk), .Q(\mem[17][19] ) );
  DFQD1 \mem_reg[17][18]  ( .D(n1524), .CP(clk), .Q(\mem[17][18] ) );
  DFQD1 \mem_reg[17][17]  ( .D(n1523), .CP(clk), .Q(\mem[17][17] ) );
  DFQD1 \mem_reg[17][16]  ( .D(n1522), .CP(clk), .Q(\mem[17][16] ) );
  DFQD1 \mem_reg[17][15]  ( .D(n1521), .CP(clk), .Q(\mem[17][15] ) );
  DFQD1 \mem_reg[17][14]  ( .D(n1520), .CP(clk), .Q(\mem[17][14] ) );
  DFQD1 \mem_reg[17][13]  ( .D(n1519), .CP(clk), .Q(\mem[17][13] ) );
  DFQD1 \mem_reg[17][12]  ( .D(n1518), .CP(clk), .Q(\mem[17][12] ) );
  DFQD1 \mem_reg[17][11]  ( .D(n1517), .CP(clk), .Q(\mem[17][11] ) );
  DFQD1 \mem_reg[17][10]  ( .D(n1516), .CP(clk), .Q(\mem[17][10] ) );
  DFQD1 \mem_reg[17][9]  ( .D(n1515), .CP(clk), .Q(\mem[17][9] ) );
  DFQD1 \mem_reg[17][8]  ( .D(n1514), .CP(clk), .Q(\mem[17][8] ) );
  DFQD1 \mem_reg[17][7]  ( .D(n1513), .CP(clk), .Q(\mem[17][7] ) );
  DFQD1 \mem_reg[17][6]  ( .D(n1512), .CP(clk), .Q(\mem[17][6] ) );
  DFQD1 \mem_reg[17][5]  ( .D(n1511), .CP(clk), .Q(\mem[17][5] ) );
  DFQD1 \mem_reg[17][4]  ( .D(n1510), .CP(clk), .Q(\mem[17][4] ) );
  DFQD1 \mem_reg[17][3]  ( .D(n1509), .CP(clk), .Q(\mem[17][3] ) );
  DFQD1 \mem_reg[17][2]  ( .D(n1508), .CP(clk), .Q(\mem[17][2] ) );
  DFQD1 \mem_reg[17][1]  ( .D(n1507), .CP(clk), .Q(\mem[17][1] ) );
  DFQD1 \mem_reg[17][0]  ( .D(n1506), .CP(clk), .Q(\mem[17][0] ) );
  DFQD1 \mem_reg[18][23]  ( .D(n1505), .CP(clk), .Q(\mem[18][23] ) );
  DFQD1 \mem_reg[18][22]  ( .D(n1504), .CP(clk), .Q(\mem[18][22] ) );
  DFQD1 \mem_reg[18][21]  ( .D(n1503), .CP(clk), .Q(\mem[18][21] ) );
  DFQD1 \mem_reg[18][20]  ( .D(n1502), .CP(clk), .Q(\mem[18][20] ) );
  DFQD1 \mem_reg[18][19]  ( .D(n1501), .CP(clk), .Q(\mem[18][19] ) );
  DFQD1 \mem_reg[18][18]  ( .D(n1500), .CP(clk), .Q(\mem[18][18] ) );
  DFQD1 \mem_reg[18][17]  ( .D(n1499), .CP(clk), .Q(\mem[18][17] ) );
  DFQD1 \mem_reg[18][16]  ( .D(n1498), .CP(clk), .Q(\mem[18][16] ) );
  DFQD1 \mem_reg[18][15]  ( .D(n1497), .CP(clk), .Q(\mem[18][15] ) );
  DFQD1 \mem_reg[18][14]  ( .D(n1496), .CP(clk), .Q(\mem[18][14] ) );
  DFQD1 \mem_reg[18][13]  ( .D(n1495), .CP(clk), .Q(\mem[18][13] ) );
  DFQD1 \mem_reg[18][12]  ( .D(n1494), .CP(clk), .Q(\mem[18][12] ) );
  DFQD1 \mem_reg[18][11]  ( .D(n1493), .CP(clk), .Q(\mem[18][11] ) );
  DFQD1 \mem_reg[18][10]  ( .D(n1492), .CP(clk), .Q(\mem[18][10] ) );
  DFQD1 \mem_reg[18][9]  ( .D(n1491), .CP(clk), .Q(\mem[18][9] ) );
  DFQD1 \mem_reg[18][8]  ( .D(n1490), .CP(clk), .Q(\mem[18][8] ) );
  DFQD1 \mem_reg[18][7]  ( .D(n1489), .CP(clk), .Q(\mem[18][7] ) );
  DFQD1 \mem_reg[18][6]  ( .D(n1488), .CP(clk), .Q(\mem[18][6] ) );
  DFQD1 \mem_reg[18][5]  ( .D(n1487), .CP(clk), .Q(\mem[18][5] ) );
  DFQD1 \mem_reg[18][4]  ( .D(n1486), .CP(clk), .Q(\mem[18][4] ) );
  DFQD1 \mem_reg[18][3]  ( .D(n1485), .CP(clk), .Q(\mem[18][3] ) );
  DFQD1 \mem_reg[18][2]  ( .D(n1484), .CP(clk), .Q(\mem[18][2] ) );
  DFQD1 \mem_reg[18][1]  ( .D(n1483), .CP(clk), .Q(\mem[18][1] ) );
  DFQD1 \mem_reg[18][0]  ( .D(n1482), .CP(clk), .Q(\mem[18][0] ) );
  DFQD1 \mem_reg[19][23]  ( .D(n1481), .CP(clk), .Q(\mem[19][23] ) );
  DFQD1 \mem_reg[19][22]  ( .D(n1480), .CP(clk), .Q(\mem[19][22] ) );
  DFQD1 \mem_reg[19][21]  ( .D(n1479), .CP(clk), .Q(\mem[19][21] ) );
  DFQD1 \mem_reg[19][20]  ( .D(n1478), .CP(clk), .Q(\mem[19][20] ) );
  DFQD1 \mem_reg[19][19]  ( .D(n1477), .CP(clk), .Q(\mem[19][19] ) );
  DFQD1 \mem_reg[19][18]  ( .D(n1476), .CP(clk), .Q(\mem[19][18] ) );
  DFQD1 \mem_reg[19][17]  ( .D(n1475), .CP(clk), .Q(\mem[19][17] ) );
  DFQD1 \mem_reg[19][16]  ( .D(n1474), .CP(clk), .Q(\mem[19][16] ) );
  DFQD1 \mem_reg[19][15]  ( .D(n1473), .CP(clk), .Q(\mem[19][15] ) );
  DFQD1 \mem_reg[19][14]  ( .D(n1472), .CP(clk), .Q(\mem[19][14] ) );
  DFQD1 \mem_reg[19][13]  ( .D(n1471), .CP(clk), .Q(\mem[19][13] ) );
  DFQD1 \mem_reg[19][12]  ( .D(n1470), .CP(clk), .Q(\mem[19][12] ) );
  DFQD1 \mem_reg[19][11]  ( .D(n1469), .CP(clk), .Q(\mem[19][11] ) );
  DFQD1 \mem_reg[19][10]  ( .D(n1468), .CP(clk), .Q(\mem[19][10] ) );
  DFQD1 \mem_reg[19][9]  ( .D(n1467), .CP(clk), .Q(\mem[19][9] ) );
  DFQD1 \mem_reg[19][8]  ( .D(n1466), .CP(clk), .Q(\mem[19][8] ) );
  DFQD1 \mem_reg[19][7]  ( .D(n1465), .CP(clk), .Q(\mem[19][7] ) );
  DFQD1 \mem_reg[19][6]  ( .D(n1464), .CP(clk), .Q(\mem[19][6] ) );
  DFQD1 \mem_reg[19][5]  ( .D(n1463), .CP(clk), .Q(\mem[19][5] ) );
  DFQD1 \mem_reg[19][4]  ( .D(n1462), .CP(clk), .Q(\mem[19][4] ) );
  DFQD1 \mem_reg[19][3]  ( .D(n1461), .CP(clk), .Q(\mem[19][3] ) );
  DFQD1 \mem_reg[19][2]  ( .D(n1460), .CP(clk), .Q(\mem[19][2] ) );
  DFQD1 \mem_reg[19][1]  ( .D(n1459), .CP(clk), .Q(\mem[19][1] ) );
  DFQD1 \mem_reg[19][0]  ( .D(n1458), .CP(clk), .Q(\mem[19][0] ) );
  DFQD1 \mem_reg[20][23]  ( .D(n1457), .CP(clk), .Q(\mem[20][23] ) );
  DFQD1 \mem_reg[20][22]  ( .D(n1456), .CP(clk), .Q(\mem[20][22] ) );
  DFQD1 \mem_reg[20][21]  ( .D(n1455), .CP(clk), .Q(\mem[20][21] ) );
  DFQD1 \mem_reg[20][20]  ( .D(n1454), .CP(clk), .Q(\mem[20][20] ) );
  DFQD1 \mem_reg[20][19]  ( .D(n1453), .CP(clk), .Q(\mem[20][19] ) );
  DFQD1 \mem_reg[20][18]  ( .D(n1452), .CP(clk), .Q(\mem[20][18] ) );
  DFQD1 \mem_reg[20][17]  ( .D(n1451), .CP(clk), .Q(\mem[20][17] ) );
  DFQD1 \mem_reg[20][16]  ( .D(n1450), .CP(clk), .Q(\mem[20][16] ) );
  DFQD1 \mem_reg[20][15]  ( .D(n1449), .CP(clk), .Q(\mem[20][15] ) );
  DFQD1 \mem_reg[20][14]  ( .D(n1448), .CP(clk), .Q(\mem[20][14] ) );
  DFQD1 \mem_reg[20][13]  ( .D(n1447), .CP(clk), .Q(\mem[20][13] ) );
  DFQD1 \mem_reg[20][12]  ( .D(n1446), .CP(clk), .Q(\mem[20][12] ) );
  DFQD1 \mem_reg[20][11]  ( .D(n1445), .CP(clk), .Q(\mem[20][11] ) );
  DFQD1 \mem_reg[20][10]  ( .D(n1444), .CP(clk), .Q(\mem[20][10] ) );
  DFQD1 \mem_reg[20][9]  ( .D(n1443), .CP(clk), .Q(\mem[20][9] ) );
  DFQD1 \mem_reg[20][8]  ( .D(n1442), .CP(clk), .Q(\mem[20][8] ) );
  DFQD1 \mem_reg[20][7]  ( .D(n1441), .CP(clk), .Q(\mem[20][7] ) );
  DFQD1 \mem_reg[20][6]  ( .D(n1440), .CP(clk), .Q(\mem[20][6] ) );
  DFQD1 \mem_reg[20][5]  ( .D(n1439), .CP(clk), .Q(\mem[20][5] ) );
  DFQD1 \mem_reg[20][4]  ( .D(n1438), .CP(clk), .Q(\mem[20][4] ) );
  DFQD1 \mem_reg[20][3]  ( .D(n1437), .CP(clk), .Q(\mem[20][3] ) );
  DFQD1 \mem_reg[20][2]  ( .D(n1436), .CP(clk), .Q(\mem[20][2] ) );
  DFQD1 \mem_reg[20][1]  ( .D(n1435), .CP(clk), .Q(\mem[20][1] ) );
  DFQD1 \mem_reg[20][0]  ( .D(n1434), .CP(clk), .Q(\mem[20][0] ) );
  DFQD1 \mem_reg[21][23]  ( .D(n1433), .CP(clk), .Q(\mem[21][23] ) );
  DFQD1 \mem_reg[21][22]  ( .D(n1432), .CP(clk), .Q(\mem[21][22] ) );
  DFQD1 \mem_reg[21][21]  ( .D(n1431), .CP(clk), .Q(\mem[21][21] ) );
  DFQD1 \mem_reg[21][20]  ( .D(n1430), .CP(clk), .Q(\mem[21][20] ) );
  DFQD1 \mem_reg[21][19]  ( .D(n1429), .CP(clk), .Q(\mem[21][19] ) );
  DFQD1 \mem_reg[21][18]  ( .D(n1428), .CP(clk), .Q(\mem[21][18] ) );
  DFQD1 \mem_reg[21][17]  ( .D(n1427), .CP(clk), .Q(\mem[21][17] ) );
  DFQD1 \mem_reg[21][16]  ( .D(n1426), .CP(clk), .Q(\mem[21][16] ) );
  DFQD1 \mem_reg[21][15]  ( .D(n1425), .CP(clk), .Q(\mem[21][15] ) );
  DFQD1 \mem_reg[21][14]  ( .D(n1424), .CP(clk), .Q(\mem[21][14] ) );
  DFQD1 \mem_reg[21][13]  ( .D(n1423), .CP(clk), .Q(\mem[21][13] ) );
  DFQD1 \mem_reg[21][12]  ( .D(n1422), .CP(clk), .Q(\mem[21][12] ) );
  DFQD1 \mem_reg[21][11]  ( .D(n1421), .CP(clk), .Q(\mem[21][11] ) );
  DFQD1 \mem_reg[21][10]  ( .D(n1420), .CP(clk), .Q(\mem[21][10] ) );
  DFQD1 \mem_reg[21][9]  ( .D(n1419), .CP(clk), .Q(\mem[21][9] ) );
  DFQD1 \mem_reg[21][8]  ( .D(n1418), .CP(clk), .Q(\mem[21][8] ) );
  DFQD1 \mem_reg[21][7]  ( .D(n1417), .CP(clk), .Q(\mem[21][7] ) );
  DFQD1 \mem_reg[21][6]  ( .D(n1416), .CP(clk), .Q(\mem[21][6] ) );
  DFQD1 \mem_reg[21][5]  ( .D(n1415), .CP(clk), .Q(\mem[21][5] ) );
  DFQD1 \mem_reg[21][4]  ( .D(n1414), .CP(clk), .Q(\mem[21][4] ) );
  DFQD1 \mem_reg[21][3]  ( .D(n1413), .CP(clk), .Q(\mem[21][3] ) );
  DFQD1 \mem_reg[21][2]  ( .D(n1412), .CP(clk), .Q(\mem[21][2] ) );
  DFQD1 \mem_reg[21][1]  ( .D(n1411), .CP(clk), .Q(\mem[21][1] ) );
  DFQD1 \mem_reg[21][0]  ( .D(n1410), .CP(clk), .Q(\mem[21][0] ) );
  DFQD1 \mem_reg[22][23]  ( .D(n1409), .CP(clk), .Q(\mem[22][23] ) );
  DFQD1 \mem_reg[22][22]  ( .D(n1408), .CP(clk), .Q(\mem[22][22] ) );
  DFQD1 \mem_reg[22][21]  ( .D(n1407), .CP(clk), .Q(\mem[22][21] ) );
  DFQD1 \mem_reg[22][20]  ( .D(n1406), .CP(clk), .Q(\mem[22][20] ) );
  DFQD1 \mem_reg[22][19]  ( .D(n1405), .CP(clk), .Q(\mem[22][19] ) );
  DFQD1 \mem_reg[22][18]  ( .D(n1404), .CP(clk), .Q(\mem[22][18] ) );
  DFQD1 \mem_reg[22][17]  ( .D(n1403), .CP(clk), .Q(\mem[22][17] ) );
  DFQD1 \mem_reg[22][16]  ( .D(n1402), .CP(clk), .Q(\mem[22][16] ) );
  DFQD1 \mem_reg[22][15]  ( .D(n1401), .CP(clk), .Q(\mem[22][15] ) );
  DFQD1 \mem_reg[22][14]  ( .D(n1400), .CP(clk), .Q(\mem[22][14] ) );
  DFQD1 \mem_reg[22][13]  ( .D(n1399), .CP(clk), .Q(\mem[22][13] ) );
  DFQD1 \mem_reg[22][12]  ( .D(n1398), .CP(clk), .Q(\mem[22][12] ) );
  DFQD1 \mem_reg[22][11]  ( .D(n1397), .CP(clk), .Q(\mem[22][11] ) );
  DFQD1 \mem_reg[22][10]  ( .D(n1396), .CP(clk), .Q(\mem[22][10] ) );
  DFQD1 \mem_reg[22][9]  ( .D(n1395), .CP(clk), .Q(\mem[22][9] ) );
  DFQD1 \mem_reg[22][8]  ( .D(n1394), .CP(clk), .Q(\mem[22][8] ) );
  DFQD1 \mem_reg[22][7]  ( .D(n1393), .CP(clk), .Q(\mem[22][7] ) );
  DFQD1 \mem_reg[22][6]  ( .D(n1392), .CP(clk), .Q(\mem[22][6] ) );
  DFQD1 \mem_reg[22][5]  ( .D(n1391), .CP(clk), .Q(\mem[22][5] ) );
  DFQD1 \mem_reg[22][4]  ( .D(n1390), .CP(clk), .Q(\mem[22][4] ) );
  DFQD1 \mem_reg[22][3]  ( .D(n1389), .CP(clk), .Q(\mem[22][3] ) );
  DFQD1 \mem_reg[22][2]  ( .D(n1388), .CP(clk), .Q(\mem[22][2] ) );
  DFQD1 \mem_reg[22][1]  ( .D(n1387), .CP(clk), .Q(\mem[22][1] ) );
  DFQD1 \mem_reg[22][0]  ( .D(n1386), .CP(clk), .Q(\mem[22][0] ) );
  DFQD1 \mem_reg[23][23]  ( .D(n1385), .CP(clk), .Q(\mem[23][23] ) );
  DFQD1 \mem_reg[23][22]  ( .D(n1384), .CP(clk), .Q(\mem[23][22] ) );
  DFQD1 \mem_reg[23][21]  ( .D(n1383), .CP(clk), .Q(\mem[23][21] ) );
  DFQD1 \mem_reg[23][20]  ( .D(n1382), .CP(clk), .Q(\mem[23][20] ) );
  DFQD1 \mem_reg[23][19]  ( .D(n1381), .CP(clk), .Q(\mem[23][19] ) );
  DFQD1 \mem_reg[23][18]  ( .D(n1380), .CP(clk), .Q(\mem[23][18] ) );
  DFQD1 \mem_reg[23][17]  ( .D(n1379), .CP(clk), .Q(\mem[23][17] ) );
  DFQD1 \mem_reg[23][16]  ( .D(n1378), .CP(clk), .Q(\mem[23][16] ) );
  DFQD1 \mem_reg[23][15]  ( .D(n1377), .CP(clk), .Q(\mem[23][15] ) );
  DFQD1 \mem_reg[23][14]  ( .D(n1376), .CP(clk), .Q(\mem[23][14] ) );
  DFQD1 \mem_reg[23][13]  ( .D(n1375), .CP(clk), .Q(\mem[23][13] ) );
  DFQD1 \mem_reg[23][12]  ( .D(n1374), .CP(clk), .Q(\mem[23][12] ) );
  DFQD1 \mem_reg[23][11]  ( .D(n1373), .CP(clk), .Q(\mem[23][11] ) );
  DFQD1 \mem_reg[23][10]  ( .D(n1372), .CP(clk), .Q(\mem[23][10] ) );
  DFQD1 \mem_reg[23][9]  ( .D(n1371), .CP(clk), .Q(\mem[23][9] ) );
  DFQD1 \mem_reg[23][8]  ( .D(n1370), .CP(clk), .Q(\mem[23][8] ) );
  DFQD1 \mem_reg[23][7]  ( .D(n1369), .CP(clk), .Q(\mem[23][7] ) );
  DFQD1 \mem_reg[23][6]  ( .D(n1368), .CP(clk), .Q(\mem[23][6] ) );
  DFQD1 \mem_reg[23][5]  ( .D(n1367), .CP(clk), .Q(\mem[23][5] ) );
  DFQD1 \mem_reg[23][4]  ( .D(n1366), .CP(clk), .Q(\mem[23][4] ) );
  DFQD1 \mem_reg[23][3]  ( .D(n1365), .CP(clk), .Q(\mem[23][3] ) );
  DFQD1 \mem_reg[23][2]  ( .D(n1364), .CP(clk), .Q(\mem[23][2] ) );
  DFQD1 \mem_reg[23][1]  ( .D(n1363), .CP(clk), .Q(\mem[23][1] ) );
  DFQD1 \mem_reg[23][0]  ( .D(n1362), .CP(clk), .Q(\mem[23][0] ) );
  DFQD1 \mem_reg[24][23]  ( .D(n1361), .CP(clk), .Q(\mem[24][23] ) );
  DFQD1 \mem_reg[24][22]  ( .D(n1360), .CP(clk), .Q(\mem[24][22] ) );
  DFQD1 \mem_reg[24][21]  ( .D(n1359), .CP(clk), .Q(\mem[24][21] ) );
  DFQD1 \mem_reg[24][20]  ( .D(n1358), .CP(clk), .Q(\mem[24][20] ) );
  DFQD1 \mem_reg[24][19]  ( .D(n1357), .CP(clk), .Q(\mem[24][19] ) );
  DFQD1 \mem_reg[24][18]  ( .D(n1356), .CP(clk), .Q(\mem[24][18] ) );
  DFQD1 \mem_reg[24][17]  ( .D(n1355), .CP(clk), .Q(\mem[24][17] ) );
  DFQD1 \mem_reg[24][16]  ( .D(n1354), .CP(clk), .Q(\mem[24][16] ) );
  DFQD1 \mem_reg[24][15]  ( .D(n1353), .CP(clk), .Q(\mem[24][15] ) );
  DFQD1 \mem_reg[24][14]  ( .D(n1352), .CP(clk), .Q(\mem[24][14] ) );
  DFQD1 \mem_reg[24][13]  ( .D(n1351), .CP(clk), .Q(\mem[24][13] ) );
  DFQD1 \mem_reg[24][12]  ( .D(n1350), .CP(clk), .Q(\mem[24][12] ) );
  DFQD1 \mem_reg[24][11]  ( .D(n1349), .CP(clk), .Q(\mem[24][11] ) );
  DFQD1 \mem_reg[24][10]  ( .D(n1348), .CP(clk), .Q(\mem[24][10] ) );
  DFQD1 \mem_reg[24][9]  ( .D(n1347), .CP(clk), .Q(\mem[24][9] ) );
  DFQD1 \mem_reg[24][8]  ( .D(n1346), .CP(clk), .Q(\mem[24][8] ) );
  DFQD1 \mem_reg[24][7]  ( .D(n1345), .CP(clk), .Q(\mem[24][7] ) );
  DFQD1 \mem_reg[24][6]  ( .D(n1344), .CP(clk), .Q(\mem[24][6] ) );
  DFQD1 \mem_reg[24][5]  ( .D(n1343), .CP(clk), .Q(\mem[24][5] ) );
  DFQD1 \mem_reg[24][4]  ( .D(n1342), .CP(clk), .Q(\mem[24][4] ) );
  DFQD1 \mem_reg[24][3]  ( .D(n1341), .CP(clk), .Q(\mem[24][3] ) );
  DFQD1 \mem_reg[24][2]  ( .D(n1340), .CP(clk), .Q(\mem[24][2] ) );
  DFQD1 \mem_reg[24][1]  ( .D(n1339), .CP(clk), .Q(\mem[24][1] ) );
  DFQD1 \mem_reg[24][0]  ( .D(n1338), .CP(clk), .Q(\mem[24][0] ) );
  DFQD1 \mem_reg[25][23]  ( .D(n1337), .CP(clk), .Q(\mem[25][23] ) );
  DFQD1 \mem_reg[25][22]  ( .D(n1336), .CP(clk), .Q(\mem[25][22] ) );
  DFQD1 \mem_reg[25][21]  ( .D(n1335), .CP(clk), .Q(\mem[25][21] ) );
  DFQD1 \mem_reg[25][20]  ( .D(n1334), .CP(clk), .Q(\mem[25][20] ) );
  DFQD1 \mem_reg[25][19]  ( .D(n1333), .CP(clk), .Q(\mem[25][19] ) );
  DFQD1 \mem_reg[25][18]  ( .D(n1332), .CP(clk), .Q(\mem[25][18] ) );
  DFQD1 \mem_reg[25][17]  ( .D(n1331), .CP(clk), .Q(\mem[25][17] ) );
  DFQD1 \mem_reg[25][16]  ( .D(n1330), .CP(clk), .Q(\mem[25][16] ) );
  DFQD1 \mem_reg[25][15]  ( .D(n1329), .CP(clk), .Q(\mem[25][15] ) );
  DFQD1 \mem_reg[25][14]  ( .D(n1328), .CP(clk), .Q(\mem[25][14] ) );
  DFQD1 \mem_reg[25][13]  ( .D(n1327), .CP(clk), .Q(\mem[25][13] ) );
  DFQD1 \mem_reg[25][12]  ( .D(n1326), .CP(clk), .Q(\mem[25][12] ) );
  DFQD1 \mem_reg[25][11]  ( .D(n1325), .CP(clk), .Q(\mem[25][11] ) );
  DFQD1 \mem_reg[25][10]  ( .D(n1324), .CP(clk), .Q(\mem[25][10] ) );
  DFQD1 \mem_reg[25][9]  ( .D(n1323), .CP(clk), .Q(\mem[25][9] ) );
  DFQD1 \mem_reg[25][8]  ( .D(n1322), .CP(clk), .Q(\mem[25][8] ) );
  DFQD1 \mem_reg[25][7]  ( .D(n1321), .CP(clk), .Q(\mem[25][7] ) );
  DFQD1 \mem_reg[25][6]  ( .D(n1320), .CP(clk), .Q(\mem[25][6] ) );
  DFQD1 \mem_reg[25][5]  ( .D(n1319), .CP(clk), .Q(\mem[25][5] ) );
  DFQD1 \mem_reg[25][4]  ( .D(n1318), .CP(clk), .Q(\mem[25][4] ) );
  DFQD1 \mem_reg[25][3]  ( .D(n1317), .CP(clk), .Q(\mem[25][3] ) );
  DFQD1 \mem_reg[25][2]  ( .D(n1316), .CP(clk), .Q(\mem[25][2] ) );
  DFQD1 \mem_reg[25][1]  ( .D(n1315), .CP(clk), .Q(\mem[25][1] ) );
  DFQD1 \mem_reg[25][0]  ( .D(n1314), .CP(clk), .Q(\mem[25][0] ) );
  DFQD1 \mem_reg[26][23]  ( .D(n1313), .CP(clk), .Q(\mem[26][23] ) );
  DFQD1 \mem_reg[26][22]  ( .D(n1312), .CP(clk), .Q(\mem[26][22] ) );
  DFQD1 \mem_reg[26][21]  ( .D(n1311), .CP(clk), .Q(\mem[26][21] ) );
  DFQD1 \mem_reg[26][20]  ( .D(n1310), .CP(clk), .Q(\mem[26][20] ) );
  DFQD1 \mem_reg[26][19]  ( .D(n1309), .CP(clk), .Q(\mem[26][19] ) );
  DFQD1 \mem_reg[26][18]  ( .D(n1308), .CP(clk), .Q(\mem[26][18] ) );
  DFQD1 \mem_reg[26][17]  ( .D(n1307), .CP(clk), .Q(\mem[26][17] ) );
  DFQD1 \mem_reg[26][16]  ( .D(n1306), .CP(clk), .Q(\mem[26][16] ) );
  DFQD1 \mem_reg[26][15]  ( .D(n1305), .CP(clk), .Q(\mem[26][15] ) );
  DFQD1 \mem_reg[26][14]  ( .D(n1304), .CP(clk), .Q(\mem[26][14] ) );
  DFQD1 \mem_reg[26][13]  ( .D(n1303), .CP(clk), .Q(\mem[26][13] ) );
  DFQD1 \mem_reg[26][12]  ( .D(n1302), .CP(clk), .Q(\mem[26][12] ) );
  DFQD1 \mem_reg[26][11]  ( .D(n1301), .CP(clk), .Q(\mem[26][11] ) );
  DFQD1 \mem_reg[26][10]  ( .D(n1300), .CP(clk), .Q(\mem[26][10] ) );
  DFQD1 \mem_reg[26][9]  ( .D(n1299), .CP(clk), .Q(\mem[26][9] ) );
  DFQD1 \mem_reg[26][8]  ( .D(n1298), .CP(clk), .Q(\mem[26][8] ) );
  DFQD1 \mem_reg[26][7]  ( .D(n1297), .CP(clk), .Q(\mem[26][7] ) );
  DFQD1 \mem_reg[26][6]  ( .D(n1296), .CP(clk), .Q(\mem[26][6] ) );
  DFQD1 \mem_reg[26][5]  ( .D(n1295), .CP(clk), .Q(\mem[26][5] ) );
  DFQD1 \mem_reg[26][4]  ( .D(n1294), .CP(clk), .Q(\mem[26][4] ) );
  DFQD1 \mem_reg[26][3]  ( .D(n1293), .CP(clk), .Q(\mem[26][3] ) );
  DFQD1 \mem_reg[26][2]  ( .D(n1292), .CP(clk), .Q(\mem[26][2] ) );
  DFQD1 \mem_reg[26][1]  ( .D(n1291), .CP(clk), .Q(\mem[26][1] ) );
  DFQD1 \mem_reg[26][0]  ( .D(n1290), .CP(clk), .Q(\mem[26][0] ) );
  DFQD1 \mem_reg[27][23]  ( .D(n1289), .CP(clk), .Q(\mem[27][23] ) );
  DFQD1 \mem_reg[27][22]  ( .D(n1288), .CP(clk), .Q(\mem[27][22] ) );
  DFQD1 \mem_reg[27][21]  ( .D(n1287), .CP(clk), .Q(\mem[27][21] ) );
  DFQD1 \mem_reg[27][20]  ( .D(n1286), .CP(clk), .Q(\mem[27][20] ) );
  DFQD1 \mem_reg[27][19]  ( .D(n1285), .CP(clk), .Q(\mem[27][19] ) );
  DFQD1 \mem_reg[27][18]  ( .D(n1284), .CP(clk), .Q(\mem[27][18] ) );
  DFQD1 \mem_reg[27][17]  ( .D(n1283), .CP(clk), .Q(\mem[27][17] ) );
  DFQD1 \mem_reg[27][16]  ( .D(n1282), .CP(clk), .Q(\mem[27][16] ) );
  DFQD1 \mem_reg[27][15]  ( .D(n1281), .CP(clk), .Q(\mem[27][15] ) );
  DFQD1 \mem_reg[27][14]  ( .D(n1280), .CP(clk), .Q(\mem[27][14] ) );
  DFQD1 \mem_reg[27][13]  ( .D(n1279), .CP(clk), .Q(\mem[27][13] ) );
  DFQD1 \mem_reg[27][12]  ( .D(n1278), .CP(clk), .Q(\mem[27][12] ) );
  DFQD1 \mem_reg[27][11]  ( .D(n1277), .CP(clk), .Q(\mem[27][11] ) );
  DFQD1 \mem_reg[27][10]  ( .D(n1276), .CP(clk), .Q(\mem[27][10] ) );
  DFQD1 \mem_reg[27][9]  ( .D(n1275), .CP(clk), .Q(\mem[27][9] ) );
  DFQD1 \mem_reg[27][8]  ( .D(n1274), .CP(clk), .Q(\mem[27][8] ) );
  DFQD1 \mem_reg[27][7]  ( .D(n1273), .CP(clk), .Q(\mem[27][7] ) );
  DFQD1 \mem_reg[27][6]  ( .D(n1272), .CP(clk), .Q(\mem[27][6] ) );
  DFQD1 \mem_reg[27][5]  ( .D(n1271), .CP(clk), .Q(\mem[27][5] ) );
  DFQD1 \mem_reg[27][4]  ( .D(n1270), .CP(clk), .Q(\mem[27][4] ) );
  DFQD1 \mem_reg[27][3]  ( .D(n1269), .CP(clk), .Q(\mem[27][3] ) );
  DFQD1 \mem_reg[27][2]  ( .D(n1268), .CP(clk), .Q(\mem[27][2] ) );
  DFQD1 \mem_reg[27][1]  ( .D(n1267), .CP(clk), .Q(\mem[27][1] ) );
  DFQD1 \mem_reg[27][0]  ( .D(n1266), .CP(clk), .Q(\mem[27][0] ) );
  DFQD1 \mem_reg[28][23]  ( .D(n1265), .CP(clk), .Q(\mem[28][23] ) );
  DFQD1 \mem_reg[28][22]  ( .D(n1264), .CP(clk), .Q(\mem[28][22] ) );
  DFQD1 \mem_reg[28][21]  ( .D(n1263), .CP(clk), .Q(\mem[28][21] ) );
  DFQD1 \mem_reg[28][20]  ( .D(n1262), .CP(clk), .Q(\mem[28][20] ) );
  DFQD1 \mem_reg[28][19]  ( .D(n1261), .CP(clk), .Q(\mem[28][19] ) );
  DFQD1 \mem_reg[28][18]  ( .D(n1260), .CP(clk), .Q(\mem[28][18] ) );
  DFQD1 \mem_reg[28][17]  ( .D(n1259), .CP(clk), .Q(\mem[28][17] ) );
  DFQD1 \mem_reg[28][16]  ( .D(n1258), .CP(clk), .Q(\mem[28][16] ) );
  DFQD1 \mem_reg[28][15]  ( .D(n1257), .CP(clk), .Q(\mem[28][15] ) );
  DFQD1 \mem_reg[28][14]  ( .D(n1256), .CP(clk), .Q(\mem[28][14] ) );
  DFQD1 \mem_reg[28][13]  ( .D(n1255), .CP(clk), .Q(\mem[28][13] ) );
  DFQD1 \mem_reg[28][12]  ( .D(n1254), .CP(clk), .Q(\mem[28][12] ) );
  DFQD1 \mem_reg[28][11]  ( .D(n1253), .CP(clk), .Q(\mem[28][11] ) );
  DFQD1 \mem_reg[28][10]  ( .D(n1252), .CP(clk), .Q(\mem[28][10] ) );
  DFQD1 \mem_reg[28][9]  ( .D(n1251), .CP(clk), .Q(\mem[28][9] ) );
  DFQD1 \mem_reg[28][8]  ( .D(n1250), .CP(clk), .Q(\mem[28][8] ) );
  DFQD1 \mem_reg[28][7]  ( .D(n1249), .CP(clk), .Q(\mem[28][7] ) );
  DFQD1 \mem_reg[28][6]  ( .D(n1248), .CP(clk), .Q(\mem[28][6] ) );
  DFQD1 \mem_reg[28][5]  ( .D(n1247), .CP(clk), .Q(\mem[28][5] ) );
  DFQD1 \mem_reg[28][4]  ( .D(n1246), .CP(clk), .Q(\mem[28][4] ) );
  DFQD1 \mem_reg[28][3]  ( .D(n1245), .CP(clk), .Q(\mem[28][3] ) );
  DFQD1 \mem_reg[28][2]  ( .D(n1244), .CP(clk), .Q(\mem[28][2] ) );
  DFQD1 \mem_reg[28][1]  ( .D(n1243), .CP(clk), .Q(\mem[28][1] ) );
  DFQD1 \mem_reg[28][0]  ( .D(n1242), .CP(clk), .Q(\mem[28][0] ) );
  DFQD1 \mem_reg[29][23]  ( .D(n1241), .CP(clk), .Q(\mem[29][23] ) );
  DFQD1 \mem_reg[29][22]  ( .D(n1240), .CP(clk), .Q(\mem[29][22] ) );
  DFQD1 \mem_reg[29][21]  ( .D(n1239), .CP(clk), .Q(\mem[29][21] ) );
  DFQD1 \mem_reg[29][20]  ( .D(n1238), .CP(clk), .Q(\mem[29][20] ) );
  DFQD1 \mem_reg[29][19]  ( .D(n1237), .CP(clk), .Q(\mem[29][19] ) );
  DFQD1 \mem_reg[29][18]  ( .D(n1236), .CP(clk), .Q(\mem[29][18] ) );
  DFQD1 \mem_reg[29][17]  ( .D(n1235), .CP(clk), .Q(\mem[29][17] ) );
  DFQD1 \mem_reg[29][16]  ( .D(n1234), .CP(clk), .Q(\mem[29][16] ) );
  DFQD1 \mem_reg[29][15]  ( .D(n1233), .CP(clk), .Q(\mem[29][15] ) );
  DFQD1 \mem_reg[29][14]  ( .D(n1232), .CP(clk), .Q(\mem[29][14] ) );
  DFQD1 \mem_reg[29][13]  ( .D(n1231), .CP(clk), .Q(\mem[29][13] ) );
  DFQD1 \mem_reg[29][12]  ( .D(n1230), .CP(clk), .Q(\mem[29][12] ) );
  DFQD1 \mem_reg[29][11]  ( .D(n1229), .CP(clk), .Q(\mem[29][11] ) );
  DFQD1 \mem_reg[29][10]  ( .D(n1228), .CP(clk), .Q(\mem[29][10] ) );
  DFQD1 \mem_reg[29][9]  ( .D(n1227), .CP(clk), .Q(\mem[29][9] ) );
  DFQD1 \mem_reg[29][8]  ( .D(n1226), .CP(clk), .Q(\mem[29][8] ) );
  DFQD1 \mem_reg[29][7]  ( .D(n1225), .CP(clk), .Q(\mem[29][7] ) );
  DFQD1 \mem_reg[29][6]  ( .D(n1224), .CP(clk), .Q(\mem[29][6] ) );
  DFQD1 \mem_reg[29][5]  ( .D(n1223), .CP(clk), .Q(\mem[29][5] ) );
  DFQD1 \mem_reg[29][4]  ( .D(n1222), .CP(clk), .Q(\mem[29][4] ) );
  DFQD1 \mem_reg[29][3]  ( .D(n1221), .CP(clk), .Q(\mem[29][3] ) );
  DFQD1 \mem_reg[29][2]  ( .D(n1220), .CP(clk), .Q(\mem[29][2] ) );
  DFQD1 \mem_reg[29][1]  ( .D(n1219), .CP(clk), .Q(\mem[29][1] ) );
  DFQD1 \mem_reg[29][0]  ( .D(n1218), .CP(clk), .Q(\mem[29][0] ) );
  DFQD1 \mem_reg[30][23]  ( .D(n1217), .CP(clk), .Q(\mem[30][23] ) );
  DFQD1 \mem_reg[30][22]  ( .D(n1216), .CP(clk), .Q(\mem[30][22] ) );
  DFQD1 \mem_reg[30][21]  ( .D(n1215), .CP(clk), .Q(\mem[30][21] ) );
  DFQD1 \mem_reg[30][20]  ( .D(n1214), .CP(clk), .Q(\mem[30][20] ) );
  DFQD1 \mem_reg[30][19]  ( .D(n1213), .CP(clk), .Q(\mem[30][19] ) );
  DFQD1 \mem_reg[30][18]  ( .D(n1212), .CP(clk), .Q(\mem[30][18] ) );
  DFQD1 \mem_reg[30][17]  ( .D(n1211), .CP(clk), .Q(\mem[30][17] ) );
  DFQD1 \mem_reg[30][16]  ( .D(n1210), .CP(clk), .Q(\mem[30][16] ) );
  DFQD1 \mem_reg[30][15]  ( .D(n1209), .CP(clk), .Q(\mem[30][15] ) );
  DFQD1 \mem_reg[30][14]  ( .D(n1208), .CP(clk), .Q(\mem[30][14] ) );
  DFQD1 \mem_reg[30][13]  ( .D(n1207), .CP(clk), .Q(\mem[30][13] ) );
  DFQD1 \mem_reg[30][12]  ( .D(n1206), .CP(clk), .Q(\mem[30][12] ) );
  DFQD1 \mem_reg[30][11]  ( .D(n1205), .CP(clk), .Q(\mem[30][11] ) );
  DFQD1 \mem_reg[30][10]  ( .D(n1204), .CP(clk), .Q(\mem[30][10] ) );
  DFQD1 \mem_reg[30][9]  ( .D(n1203), .CP(clk), .Q(\mem[30][9] ) );
  DFQD1 \mem_reg[30][8]  ( .D(n1202), .CP(clk), .Q(\mem[30][8] ) );
  DFQD1 \mem_reg[30][7]  ( .D(n1201), .CP(clk), .Q(\mem[30][7] ) );
  DFQD1 \mem_reg[30][6]  ( .D(n1200), .CP(clk), .Q(\mem[30][6] ) );
  DFQD1 \mem_reg[30][5]  ( .D(n1199), .CP(clk), .Q(\mem[30][5] ) );
  DFQD1 \mem_reg[30][4]  ( .D(n1198), .CP(clk), .Q(\mem[30][4] ) );
  DFQD1 \mem_reg[30][3]  ( .D(n1197), .CP(clk), .Q(\mem[30][3] ) );
  DFQD1 \mem_reg[30][2]  ( .D(n1196), .CP(clk), .Q(\mem[30][2] ) );
  DFQD1 \mem_reg[30][1]  ( .D(n1195), .CP(clk), .Q(\mem[30][1] ) );
  DFQD1 \mem_reg[30][0]  ( .D(n1194), .CP(clk), .Q(\mem[30][0] ) );
  DFQD1 \mem_reg[31][23]  ( .D(n1193), .CP(clk), .Q(\mem[31][23] ) );
  DFQD1 \mem_reg[31][22]  ( .D(n1192), .CP(clk), .Q(\mem[31][22] ) );
  DFQD1 \mem_reg[31][21]  ( .D(n1191), .CP(clk), .Q(\mem[31][21] ) );
  DFQD1 \mem_reg[31][20]  ( .D(n1190), .CP(clk), .Q(\mem[31][20] ) );
  DFQD1 \mem_reg[31][19]  ( .D(n1189), .CP(clk), .Q(\mem[31][19] ) );
  DFQD1 \mem_reg[31][18]  ( .D(n1188), .CP(clk), .Q(\mem[31][18] ) );
  DFQD1 \mem_reg[31][17]  ( .D(n1187), .CP(clk), .Q(\mem[31][17] ) );
  DFQD1 \mem_reg[31][16]  ( .D(n1186), .CP(clk), .Q(\mem[31][16] ) );
  DFQD1 \mem_reg[31][15]  ( .D(n1185), .CP(clk), .Q(\mem[31][15] ) );
  DFQD1 \mem_reg[31][14]  ( .D(n1184), .CP(clk), .Q(\mem[31][14] ) );
  DFQD1 \mem_reg[31][13]  ( .D(n1183), .CP(clk), .Q(\mem[31][13] ) );
  DFQD1 \mem_reg[31][12]  ( .D(n1182), .CP(clk), .Q(\mem[31][12] ) );
  DFQD1 \mem_reg[31][11]  ( .D(n1181), .CP(clk), .Q(\mem[31][11] ) );
  DFQD1 \mem_reg[31][10]  ( .D(n1180), .CP(clk), .Q(\mem[31][10] ) );
  DFQD1 \mem_reg[31][9]  ( .D(n1179), .CP(clk), .Q(\mem[31][9] ) );
  DFQD1 \mem_reg[31][8]  ( .D(n1178), .CP(clk), .Q(\mem[31][8] ) );
  DFQD1 \mem_reg[31][7]  ( .D(n1177), .CP(clk), .Q(\mem[31][7] ) );
  DFQD1 \mem_reg[31][6]  ( .D(n1176), .CP(clk), .Q(\mem[31][6] ) );
  DFQD1 \mem_reg[31][5]  ( .D(n1175), .CP(clk), .Q(\mem[31][5] ) );
  DFQD1 \mem_reg[31][4]  ( .D(n1174), .CP(clk), .Q(\mem[31][4] ) );
  DFQD1 \mem_reg[31][3]  ( .D(n1173), .CP(clk), .Q(\mem[31][3] ) );
  DFQD1 \mem_reg[31][2]  ( .D(n1172), .CP(clk), .Q(\mem[31][2] ) );
  DFQD1 \mem_reg[31][1]  ( .D(n1171), .CP(clk), .Q(\mem[31][1] ) );
  DFQD1 \mem_reg[31][0]  ( .D(n1170), .CP(clk), .Q(\mem[31][0] ) );
  CKND2D0 U2 ( .A1(dirb[2]), .A2(n18), .ZN(n19) );
  INVD0 U3 ( .I(dira[4]), .ZN(n87) );
  NR2D0 U4 ( .A1(n9), .A2(n7), .ZN(n8) );
  CKND2D0 U5 ( .A1(dira[2]), .A2(n224), .ZN(n80) );
  AOI22D0 U6 ( .A1(\mem[24][0] ), .A2(n774), .B1(\mem[26][0] ), .B2(n773), 
        .ZN(n58) );
  AOI22D0 U7 ( .A1(n774), .A2(\mem[24][1] ), .B1(n773), .B2(\mem[26][1] ), 
        .ZN(n511) );
  AOI22D0 U8 ( .A1(n764), .A2(\mem[13][2] ), .B1(n763), .B2(\mem[15][2] ), 
        .ZN(n765) );
  AOI22D0 U9 ( .A1(n758), .A2(\mem[11][3] ), .B1(n757), .B2(\mem[4][3] ), .ZN(
        n487) );
  AOI22D0 U10 ( .A1(n784), .A2(\mem[21][5] ), .B1(n783), .B2(\mem[23][5] ), 
        .ZN(n472) );
  AOI22D0 U11 ( .A1(n774), .A2(\mem[24][6] ), .B1(n773), .B2(\mem[26][6] ), 
        .ZN(n555) );
  AOI22D0 U12 ( .A1(n764), .A2(\mem[13][7] ), .B1(n763), .B2(\mem[15][7] ), 
        .ZN(n440) );
  AOI22D0 U13 ( .A1(n758), .A2(\mem[11][8] ), .B1(n757), .B2(\mem[4][8] ), 
        .ZN(n575) );
  AOI22D0 U14 ( .A1(n784), .A2(\mem[21][10] ), .B1(n783), .B2(\mem[23][10] ), 
        .ZN(n604) );
  AOI22D0 U15 ( .A1(n774), .A2(\mem[24][11] ), .B1(n773), .B2(\mem[26][11] ), 
        .ZN(n401) );
  AOI22D0 U16 ( .A1(n764), .A2(\mem[13][12] ), .B1(n763), .B2(\mem[15][12] ), 
        .ZN(n616) );
  AOI22D0 U17 ( .A1(n758), .A2(\mem[11][13] ), .B1(n757), .B2(\mem[4][13] ), 
        .ZN(n377) );
  AOI22D0 U18 ( .A1(n784), .A2(\mem[21][15] ), .B1(n783), .B2(\mem[23][15] ), 
        .ZN(n362) );
  AOI22D0 U19 ( .A1(n774), .A2(\mem[24][16] ), .B1(n773), .B2(\mem[26][16] ), 
        .ZN(n665) );
  AOI22D0 U20 ( .A1(n764), .A2(\mem[13][17] ), .B1(n763), .B2(\mem[15][17] ), 
        .ZN(n330) );
  AOI22D0 U21 ( .A1(n758), .A2(\mem[11][18] ), .B1(n757), .B2(\mem[4][18] ), 
        .ZN(n685) );
  AOI22D0 U22 ( .A1(n784), .A2(\mem[21][20] ), .B1(n783), .B2(\mem[23][20] ), 
        .ZN(n714) );
  AOI22D0 U23 ( .A1(n774), .A2(\mem[24][21] ), .B1(n773), .B2(\mem[26][21] ), 
        .ZN(n291) );
  AOI22D0 U24 ( .A1(n764), .A2(\mem[13][22] ), .B1(n763), .B2(\mem[15][22] ), 
        .ZN(n726) );
  AOI22D0 U25 ( .A1(n758), .A2(\mem[11][23] ), .B1(n757), .B2(\mem[4][23] ), 
        .ZN(n23) );
  AOI22D0 U26 ( .A1(\mem[1][1] ), .A2(n1123), .B1(\mem[3][1] ), .B2(n1122), 
        .ZN(n1022) );
  AOI22D0 U27 ( .A1(\mem[8][2] ), .A2(n1125), .B1(\mem[10][2] ), .B2(n1124), 
        .ZN(n165) );
  AOI22D0 U28 ( .A1(\mem[11][3] ), .A2(n1127), .B1(\mem[9][3] ), .B2(n1126), 
        .ZN(n1060) );
  AOI22D0 U29 ( .A1(\mem[4][4] ), .A2(n1133), .B1(\mem[6][4] ), .B2(n1132), 
        .ZN(n1007) );
  AOI22D0 U30 ( .A1(\mem[5][5] ), .A2(n1135), .B1(\mem[7][5] ), .B2(n1134), 
        .ZN(n150) );
  AOI22D0 U31 ( .A1(\mem[12][6] ), .A2(n1137), .B1(\mem[14][6] ), .B2(n1136), 
        .ZN(n985) );
  AOI22D0 U32 ( .A1(\mem[13][7] ), .A2(n1139), .B1(\mem[15][7] ), .B2(n1138), 
        .ZN(n964) );
  AOI22D0 U33 ( .A1(\mem[16][8] ), .A2(n1145), .B1(\mem[18][8] ), .B2(n1144), 
        .ZN(n135) );
  AOI22D0 U34 ( .A1(\mem[17][9] ), .A2(n1147), .B1(\mem[19][9] ), .B2(n1146), 
        .ZN(n1090) );
  AOI22D0 U35 ( .A1(\mem[24][10] ), .A2(n1149), .B1(\mem[26][10] ), .B2(n1148), 
        .ZN(n949) );
  AOI22D0 U36 ( .A1(\mem[25][11] ), .A2(n1151), .B1(\mem[27][11] ), .B2(n1150), 
        .ZN(n192) );
  AOI22D0 U37 ( .A1(\mem[20][12] ), .A2(n1157), .B1(\mem[22][12] ), .B2(n1156), 
        .ZN(n935) );
  AOI22D0 U38 ( .A1(\mem[21][13] ), .A2(n1159), .B1(\mem[23][13] ), .B2(n1158), 
        .ZN(n914) );
  AOI22D0 U39 ( .A1(\mem[28][14] ), .A2(n1161), .B1(\mem[30][14] ), .B2(n1160), 
        .ZN(n117) );
  AOI22D0 U40 ( .A1(\mem[29][15] ), .A2(n1163), .B1(\mem[31][15] ), .B2(n1162), 
        .ZN(n1112) );
  AOI22D0 U41 ( .A1(\mem[0][15] ), .A2(n1121), .B1(\mem[2][15] ), .B2(n1120), 
        .ZN(n1103) );
  AOI22D0 U42 ( .A1(\mem[1][16] ), .A2(n1123), .B1(\mem[3][16] ), .B2(n1122), 
        .ZN(n882) );
  AOI22D0 U43 ( .A1(\mem[8][17] ), .A2(n1125), .B1(\mem[10][17] ), .B2(n1124), 
        .ZN(n205) );
  AOI22D0 U44 ( .A1(\mem[11][18] ), .A2(n1127), .B1(\mem[9][18] ), .B2(n1126), 
        .ZN(n860) );
  AOI22D0 U45 ( .A1(\mem[4][19] ), .A2(n1133), .B1(\mem[6][19] ), .B2(n1132), 
        .ZN(n847) );
  AOI22D0 U46 ( .A1(\mem[5][20] ), .A2(n1135), .B1(\mem[7][20] ), .B2(n1134), 
        .ZN(n84) );
  AOI22D0 U47 ( .A1(\mem[12][21] ), .A2(n1137), .B1(\mem[14][21] ), .B2(n1136), 
        .ZN(n1141) );
  AOI22D0 U48 ( .A1(\mem[13][22] ), .A2(n1139), .B1(\mem[15][22] ), .B2(n1138), 
        .ZN(n824) );
  AOI22D0 U49 ( .A1(\mem[16][23] ), .A2(n1145), .B1(\mem[18][23] ), .B2(n1144), 
        .ZN(n811) );
  ND4D0 U50 ( .A1(n495), .A2(n494), .A3(n493), .A4(n492), .ZN(n496) );
  ND4D0 U51 ( .A1(n561), .A2(n560), .A3(n559), .A4(n558), .ZN(n562) );
  ND4D0 U52 ( .A1(n429), .A2(n428), .A3(n427), .A4(n426), .ZN(n430) );
  ND4D0 U53 ( .A1(n627), .A2(n626), .A3(n625), .A4(n624), .ZN(n628) );
  ND4D0 U54 ( .A1(n363), .A2(n362), .A3(n361), .A4(n360), .ZN(n364) );
  ND4D0 U55 ( .A1(n693), .A2(n692), .A3(n691), .A4(n690), .ZN(n694) );
  ND4D0 U56 ( .A1(n297), .A2(n296), .A3(n295), .A4(n294), .ZN(n298) );
  INVD0 U57 ( .I(n9), .ZN(n756) );
  AOI22D0 U58 ( .A1(\mem[5][0] ), .A2(n1135), .B1(\mem[7][0] ), .B2(n1134), 
        .ZN(n1046) );
  INVD0 U59 ( .I(data[8]), .ZN(n571) );
  ND4D0 U60 ( .A1(n1035), .A2(n1034), .A3(n1033), .A4(n1032), .ZN(n1036) );
  ND4D0 U61 ( .A1(n1003), .A2(n1002), .A3(n1001), .A4(n1000), .ZN(n1019) );
  ND4D0 U62 ( .A1(n131), .A2(n130), .A3(n129), .A4(n128), .ZN(n142) );
  ND4D0 U63 ( .A1(n931), .A2(n930), .A3(n929), .A4(n928), .ZN(n937) );
  ND4D0 U64 ( .A1(n895), .A2(n894), .A3(n893), .A4(n892), .ZN(n896) );
  ND4D0 U65 ( .A1(n843), .A2(n842), .A3(n841), .A4(n840), .ZN(n859) );
  ND4D0 U66 ( .A1(n807), .A2(n806), .A3(n805), .A4(n804), .ZN(n818) );
  AOI22D0 U67 ( .A1(n746), .A2(\mem[30][2] ), .B1(n745), .B2(\mem[2][2] ), 
        .ZN(n799) );
  AOI22D0 U68 ( .A1(n748), .A2(\mem[1][6] ), .B1(n747), .B2(\mem[3][6] ), .ZN(
        n567) );
  OA211D0 U69 ( .A1(n756), .A2(n593), .B(n592), .C(n591), .Z(n610) );
  OA211D0 U70 ( .A1(n756), .A2(n637), .B(n636), .C(n635), .Z(n654) );
  AOI22D0 U71 ( .A1(n746), .A2(\mem[30][17] ), .B1(n745), .B2(\mem[2][17] ), 
        .ZN(n348) );
  AOI22D0 U72 ( .A1(n748), .A2(\mem[1][21] ), .B1(n747), .B2(\mem[3][21] ), 
        .ZN(n303) );
  MAOI22D0 U73 ( .A1(n252), .A2(n281), .B1(\mem[31][0] ), .B2(n252), .ZN(n1170) );
  MAOI22D0 U74 ( .A1(n252), .A2(n637), .B1(\mem[31][14] ), .B2(n252), .ZN(
        n1184) );
  MAOI22D0 U75 ( .A1(n253), .A2(n461), .B1(\mem[30][5] ), .B2(n253), .ZN(n1199) );
  MAOI22D0 U76 ( .A1(n253), .A2(n703), .B1(\mem[30][20] ), .B2(n253), .ZN(
        n1214) );
  MAOI22D0 U77 ( .A1(n255), .A2(n395), .B1(\mem[29][11] ), .B2(n255), .ZN(
        n1229) );
  MAOI22D0 U78 ( .A1(n256), .A2(n755), .B1(\mem[28][2] ), .B2(n256), .ZN(n1244) );
  MAOI22D0 U79 ( .A1(n256), .A2(n329), .B1(\mem[28][17] ), .B2(n256), .ZN(
        n1259) );
  MAOI22D0 U80 ( .A1(n245), .A2(n571), .B1(\mem[27][8] ), .B2(n245), .ZN(n1274) );
  MAOI22D0 U81 ( .A1(n245), .A2(n279), .B1(\mem[27][23] ), .B2(n245), .ZN(
        n1289) );
  MAOI22D0 U82 ( .A1(n246), .A2(n637), .B1(\mem[26][14] ), .B2(n246), .ZN(
        n1304) );
  MAOI22D0 U83 ( .A1(n247), .A2(n461), .B1(\mem[25][5] ), .B2(n247), .ZN(n1319) );
  MAOI22D0 U84 ( .A1(n247), .A2(n703), .B1(\mem[25][20] ), .B2(n247), .ZN(
        n1334) );
  MAOI22D0 U85 ( .A1(n248), .A2(n395), .B1(\mem[24][11] ), .B2(n248), .ZN(
        n1349) );
  MAOI22D0 U86 ( .A1(n250), .A2(n755), .B1(\mem[23][2] ), .B2(n250), .ZN(n1364) );
  MAOI22D0 U87 ( .A1(n250), .A2(n329), .B1(\mem[23][17] ), .B2(n250), .ZN(
        n1379) );
  MAOI22D0 U88 ( .A1(n251), .A2(n571), .B1(\mem[22][8] ), .B2(n251), .ZN(n1394) );
  MAOI22D0 U89 ( .A1(n251), .A2(n279), .B1(\mem[22][23] ), .B2(n251), .ZN(
        n1409) );
  MAOI22D0 U90 ( .A1(n273), .A2(n637), .B1(\mem[21][14] ), .B2(n273), .ZN(
        n1424) );
  MAOI22D0 U91 ( .A1(n269), .A2(n461), .B1(\mem[20][5] ), .B2(n269), .ZN(n1439) );
  MAOI22D0 U92 ( .A1(n269), .A2(n703), .B1(\mem[20][20] ), .B2(n269), .ZN(
        n1454) );
  MAOI22D0 U93 ( .A1(n271), .A2(n395), .B1(\mem[19][11] ), .B2(n271), .ZN(
        n1469) );
  MAOI22D0 U94 ( .A1(n274), .A2(n755), .B1(\mem[18][2] ), .B2(n274), .ZN(n1484) );
  MAOI22D0 U95 ( .A1(n274), .A2(n329), .B1(\mem[18][17] ), .B2(n274), .ZN(
        n1499) );
  MAOI22D0 U96 ( .A1(n276), .A2(n571), .B1(\mem[17][8] ), .B2(n276), .ZN(n1514) );
  MAOI22D0 U97 ( .A1(n276), .A2(n279), .B1(\mem[17][23] ), .B2(n276), .ZN(
        n1529) );
  MAOI22D0 U98 ( .A1(n280), .A2(n637), .B1(\mem[16][14] ), .B2(n280), .ZN(
        n1544) );
  MAOI22D0 U99 ( .A1(n282), .A2(n461), .B1(\mem[15][5] ), .B2(n282), .ZN(n1559) );
  MAOI22D0 U100 ( .A1(n282), .A2(n703), .B1(\mem[15][20] ), .B2(n282), .ZN(
        n1574) );
  MAOI22D0 U101 ( .A1(n259), .A2(n395), .B1(\mem[14][11] ), .B2(n259), .ZN(
        n1589) );
  MAOI22D0 U102 ( .A1(n261), .A2(n755), .B1(\mem[13][2] ), .B2(n261), .ZN(
        n1604) );
  MAOI22D0 U103 ( .A1(n261), .A2(n329), .B1(\mem[13][17] ), .B2(n261), .ZN(
        n1619) );
  MAOI22D0 U104 ( .A1(n262), .A2(n571), .B1(\mem[12][8] ), .B2(n262), .ZN(
        n1634) );
  MAOI22D0 U105 ( .A1(n262), .A2(n279), .B1(\mem[12][23] ), .B2(n262), .ZN(
        n1649) );
  MAOI22D0 U106 ( .A1(n263), .A2(n637), .B1(\mem[11][14] ), .B2(n263), .ZN(
        n1664) );
  MAOI22D0 U107 ( .A1(n264), .A2(n461), .B1(\mem[10][5] ), .B2(n264), .ZN(
        n1679) );
  MAOI22D0 U108 ( .A1(n264), .A2(n703), .B1(\mem[10][20] ), .B2(n264), .ZN(
        n1694) );
  MAOI22D0 U109 ( .A1(n266), .A2(n395), .B1(\mem[9][11] ), .B2(n266), .ZN(
        n1709) );
  MAOI22D0 U110 ( .A1(n267), .A2(n755), .B1(\mem[8][2] ), .B2(n267), .ZN(n1724) );
  MAOI22D0 U111 ( .A1(n267), .A2(n329), .B1(\mem[8][17] ), .B2(n267), .ZN(
        n1739) );
  MAOI22D0 U112 ( .A1(n231), .A2(n571), .B1(\mem[7][8] ), .B2(n231), .ZN(n1754) );
  MAOI22D0 U113 ( .A1(n231), .A2(n279), .B1(\mem[7][23] ), .B2(n231), .ZN(
        n1769) );
  MAOI22D0 U114 ( .A1(n233), .A2(n637), .B1(\mem[6][14] ), .B2(n233), .ZN(
        n1784) );
  MAOI22D0 U115 ( .A1(n235), .A2(n461), .B1(\mem[5][5] ), .B2(n235), .ZN(n1799) );
  MAOI22D0 U116 ( .A1(n235), .A2(n703), .B1(\mem[5][20] ), .B2(n235), .ZN(
        n1814) );
  MAOI22D0 U117 ( .A1(n237), .A2(n395), .B1(\mem[4][11] ), .B2(n237), .ZN(
        n1829) );
  MAOI22D0 U118 ( .A1(n239), .A2(n755), .B1(\mem[3][2] ), .B2(n239), .ZN(n1844) );
  MAOI22D0 U119 ( .A1(n239), .A2(n329), .B1(\mem[3][17] ), .B2(n239), .ZN(
        n1859) );
  MAOI22D0 U120 ( .A1(n243), .A2(n571), .B1(\mem[2][8] ), .B2(n243), .ZN(n1874) );
  MAOI22D0 U121 ( .A1(n243), .A2(n279), .B1(\mem[2][23] ), .B2(n243), .ZN(
        n1889) );
  MAOI22D0 U122 ( .A1(n228), .A2(n637), .B1(\mem[1][14] ), .B2(n228), .ZN(
        n1904) );
  MAOI22D0 U123 ( .A1(n227), .A2(n461), .B1(\mem[0][5] ), .B2(n227), .ZN(n1919) );
  MAOI22D0 U124 ( .A1(n227), .A2(n703), .B1(\mem[0][20] ), .B2(n227), .ZN(
        n1934) );
  ND4D0 U125 ( .A1(n458), .A2(n457), .A3(n456), .A4(n455), .ZN(B[7]) );
  ND4D0 U126 ( .A1(n744), .A2(n743), .A3(n742), .A4(n741), .ZN(B[22]) );
  INVD0 U127 ( .I(dira[0]), .ZN(n72) );
  INVD0 U128 ( .I(dirb[0]), .ZN(n11) );
  INVD0 U129 ( .I(dirb[3]), .ZN(n10) );
  INVD0 U130 ( .I(dirb[4]), .ZN(n13) );
  OAI22D0 U131 ( .A1(dira[4]), .A2(n13), .B1(dira[3]), .B2(n10), .ZN(n1) );
  AOI221D0 U132 ( .A1(n10), .A2(dira[3]), .B1(n13), .B2(dira[4]), .C(n1), .ZN(
        n4) );
  INVD0 U133 ( .I(dira[1]), .ZN(n73) );
  INVD0 U134 ( .I(dirb[1]), .ZN(n7) );
  INVD0 U135 ( .I(dirb[2]), .ZN(n26) );
  INVD0 U136 ( .I(dira[2]), .ZN(n240) );
  OAI221D0 U137 ( .A1(dira[2]), .A2(n26), .B1(n240), .B2(dirb[2]), .C(write), 
        .ZN(n2) );
  AOI221D0 U138 ( .A1(dirb[1]), .A2(n73), .B1(n7), .B2(dira[1]), .C(n2), .ZN(
        n3) );
  CKND2D0 U139 ( .A1(n4), .A2(n3), .ZN(n5) );
  AOI221D0 U140 ( .A1(dirb[0]), .A2(n72), .B1(n11), .B2(dira[0]), .C(n5), .ZN(
        n9) );
  NR2D0 U141 ( .A1(dirb[0]), .A2(n9), .ZN(n6) );
  CKND2D0 U142 ( .A1(dirb[1]), .A2(n6), .ZN(n33) );
  ND3D0 U143 ( .A1(dirb[2]), .A2(dirb[3]), .A3(dirb[4]), .ZN(n36) );
  NR2D0 U144 ( .A1(n33), .A2(n36), .ZN(n746) );
  NR2D0 U145 ( .A1(dirb[2]), .A2(dirb[3]), .ZN(n24) );
  CKND2D0 U146 ( .A1(n24), .A2(n13), .ZN(n38) );
  NR2D0 U147 ( .A1(n33), .A2(n38), .ZN(n745) );
  AOI22D0 U148 ( .A1(n746), .A2(\mem[30][23] ), .B1(n745), .B2(\mem[2][23] ), 
        .ZN(n50) );
  NR2D0 U149 ( .A1(dirb[1]), .A2(n9), .ZN(n12) );
  CKND2D0 U150 ( .A1(dirb[0]), .A2(n12), .ZN(n35) );
  NR2D0 U151 ( .A1(n35), .A2(n38), .ZN(n748) );
  CKND2D0 U152 ( .A1(dirb[0]), .A2(n8), .ZN(n37) );
  NR2D0 U153 ( .A1(n37), .A2(n38), .ZN(n747) );
  AOI22D0 U154 ( .A1(n748), .A2(\mem[1][23] ), .B1(n747), .B2(\mem[3][23] ), 
        .ZN(n49) );
  INVD0 U155 ( .I(data[23]), .ZN(n279) );
  NR2D0 U156 ( .A1(dirb[4]), .A2(n10), .ZN(n18) );
  CKND2D0 U157 ( .A1(n18), .A2(n26), .ZN(n16) );
  CKND2D0 U158 ( .A1(n12), .A2(n11), .ZN(n39) );
  NR2D0 U159 ( .A1(n16), .A2(n39), .ZN(n750) );
  NR2D0 U160 ( .A1(n16), .A2(n33), .ZN(n749) );
  AOI22D0 U161 ( .A1(n750), .A2(\mem[8][23] ), .B1(n749), .B2(\mem[10][23] ), 
        .ZN(n15) );
  NR2D0 U162 ( .A1(dirb[3]), .A2(n26), .ZN(n32) );
  CKND2D0 U163 ( .A1(n32), .A2(n13), .ZN(n17) );
  NR2D0 U164 ( .A1(n17), .A2(n33), .ZN(n752) );
  NR2D0 U165 ( .A1(n16), .A2(n35), .ZN(n751) );
  AOI22D0 U166 ( .A1(n752), .A2(\mem[6][23] ), .B1(n751), .B2(\mem[9][23] ), 
        .ZN(n14) );
  OA211D0 U167 ( .A1(n756), .A2(n279), .B(n15), .C(n14), .Z(n48) );
  NR2D0 U168 ( .A1(n37), .A2(n16), .ZN(n758) );
  NR2D0 U169 ( .A1(n17), .A2(n39), .ZN(n757) );
  NR2D0 U170 ( .A1(n17), .A2(n35), .ZN(n760) );
  NR2D0 U171 ( .A1(n37), .A2(n17), .ZN(n759) );
  AOI22D0 U172 ( .A1(n760), .A2(\mem[5][23] ), .B1(n759), .B2(\mem[7][23] ), 
        .ZN(n22) );
  NR2D0 U173 ( .A1(n39), .A2(n19), .ZN(n762) );
  NR2D0 U174 ( .A1(n19), .A2(n33), .ZN(n761) );
  AOI22D0 U175 ( .A1(n762), .A2(\mem[12][23] ), .B1(n761), .B2(\mem[14][23] ), 
        .ZN(n21) );
  NR2D0 U176 ( .A1(n35), .A2(n19), .ZN(n764) );
  NR2D0 U177 ( .A1(n37), .A2(n19), .ZN(n763) );
  AOI22D0 U178 ( .A1(n764), .A2(\mem[13][23] ), .B1(n763), .B2(\mem[15][23] ), 
        .ZN(n20) );
  ND4D0 U179 ( .A1(n23), .A2(n22), .A3(n21), .A4(n20), .ZN(n46) );
  CKND2D0 U180 ( .A1(dirb[4]), .A2(n24), .ZN(n25) );
  NR2D0 U181 ( .A1(n39), .A2(n25), .ZN(n770) );
  NR2D0 U182 ( .A1(n33), .A2(n25), .ZN(n769) );
  AOI22D0 U183 ( .A1(n770), .A2(\mem[16][23] ), .B1(n769), .B2(\mem[18][23] ), 
        .ZN(n31) );
  NR2D0 U184 ( .A1(n35), .A2(n25), .ZN(n772) );
  NR2D0 U185 ( .A1(n37), .A2(n25), .ZN(n771) );
  AOI22D0 U186 ( .A1(n772), .A2(\mem[17][23] ), .B1(n771), .B2(\mem[19][23] ), 
        .ZN(n30) );
  ND3D0 U187 ( .A1(dirb[3]), .A2(dirb[4]), .A3(n26), .ZN(n27) );
  NR2D0 U188 ( .A1(n39), .A2(n27), .ZN(n774) );
  NR2D0 U189 ( .A1(n33), .A2(n27), .ZN(n773) );
  AOI22D0 U190 ( .A1(n774), .A2(\mem[24][23] ), .B1(n773), .B2(\mem[26][23] ), 
        .ZN(n29) );
  NR2D0 U191 ( .A1(n35), .A2(n27), .ZN(n776) );
  NR2D0 U192 ( .A1(n37), .A2(n27), .ZN(n775) );
  AOI22D0 U193 ( .A1(n776), .A2(\mem[25][23] ), .B1(n775), .B2(\mem[27][23] ), 
        .ZN(n28) );
  ND4D0 U194 ( .A1(n31), .A2(n30), .A3(n29), .A4(n28), .ZN(n45) );
  CKND2D0 U195 ( .A1(dirb[4]), .A2(n32), .ZN(n34) );
  NR2D0 U196 ( .A1(n39), .A2(n34), .ZN(n782) );
  NR2D0 U197 ( .A1(n33), .A2(n34), .ZN(n781) );
  AOI22D0 U198 ( .A1(n782), .A2(\mem[20][23] ), .B1(n781), .B2(\mem[22][23] ), 
        .ZN(n43) );
  NR2D0 U199 ( .A1(n35), .A2(n34), .ZN(n784) );
  NR2D0 U200 ( .A1(n37), .A2(n34), .ZN(n783) );
  AOI22D0 U201 ( .A1(n784), .A2(\mem[21][23] ), .B1(n783), .B2(\mem[23][23] ), 
        .ZN(n42) );
  NR2D0 U202 ( .A1(n39), .A2(n36), .ZN(n786) );
  NR2D0 U203 ( .A1(n35), .A2(n36), .ZN(n785) );
  AOI22D0 U204 ( .A1(n786), .A2(\mem[28][23] ), .B1(n785), .B2(\mem[29][23] ), 
        .ZN(n41) );
  NR2D0 U205 ( .A1(n37), .A2(n36), .ZN(n788) );
  NR2D0 U206 ( .A1(n39), .A2(n38), .ZN(n787) );
  AOI22D0 U207 ( .A1(n788), .A2(\mem[31][23] ), .B1(n787), .B2(\mem[0][23] ), 
        .ZN(n40) );
  ND4D0 U208 ( .A1(n43), .A2(n42), .A3(n41), .A4(n40), .ZN(n44) );
  NR3D0 U209 ( .A1(n46), .A2(n45), .A3(n44), .ZN(n47) );
  ND4D0 U210 ( .A1(n50), .A2(n49), .A3(n48), .A4(n47), .ZN(B[23]) );
  AOI22D0 U211 ( .A1(\mem[30][0] ), .A2(n746), .B1(\mem[2][0] ), .B2(n745), 
        .ZN(n71) );
  AOI22D0 U212 ( .A1(\mem[1][0] ), .A2(n748), .B1(\mem[3][0] ), .B2(n747), 
        .ZN(n70) );
  INVD0 U213 ( .I(data[0]), .ZN(n281) );
  AOI22D0 U214 ( .A1(\mem[8][0] ), .A2(n750), .B1(\mem[10][0] ), .B2(n749), 
        .ZN(n52) );
  AOI22D0 U215 ( .A1(\mem[6][0] ), .A2(n752), .B1(\mem[9][0] ), .B2(n751), 
        .ZN(n51) );
  OA211D0 U216 ( .A1(n756), .A2(n281), .B(n52), .C(n51), .Z(n69) );
  AOI22D0 U217 ( .A1(\mem[11][0] ), .A2(n758), .B1(\mem[4][0] ), .B2(n757), 
        .ZN(n56) );
  AOI22D0 U218 ( .A1(\mem[5][0] ), .A2(n760), .B1(\mem[7][0] ), .B2(n759), 
        .ZN(n55) );
  AOI22D0 U219 ( .A1(\mem[12][0] ), .A2(n762), .B1(\mem[14][0] ), .B2(n761), 
        .ZN(n54) );
  AOI22D0 U220 ( .A1(\mem[13][0] ), .A2(n764), .B1(\mem[15][0] ), .B2(n763), 
        .ZN(n53) );
  ND4D0 U221 ( .A1(n56), .A2(n55), .A3(n54), .A4(n53), .ZN(n67) );
  AOI22D0 U222 ( .A1(\mem[16][0] ), .A2(n770), .B1(\mem[18][0] ), .B2(n769), 
        .ZN(n60) );
  AOI22D0 U223 ( .A1(\mem[17][0] ), .A2(n772), .B1(\mem[19][0] ), .B2(n771), 
        .ZN(n59) );
  AOI22D0 U224 ( .A1(\mem[25][0] ), .A2(n776), .B1(\mem[27][0] ), .B2(n775), 
        .ZN(n57) );
  ND4D0 U225 ( .A1(n60), .A2(n59), .A3(n58), .A4(n57), .ZN(n66) );
  AOI22D0 U226 ( .A1(\mem[20][0] ), .A2(n782), .B1(\mem[22][0] ), .B2(n781), 
        .ZN(n64) );
  AOI22D0 U227 ( .A1(\mem[21][0] ), .A2(n784), .B1(\mem[23][0] ), .B2(n783), 
        .ZN(n63) );
  AOI22D0 U228 ( .A1(\mem[28][0] ), .A2(n786), .B1(\mem[29][0] ), .B2(n785), 
        .ZN(n62) );
  AOI22D0 U229 ( .A1(\mem[31][0] ), .A2(n788), .B1(\mem[0][0] ), .B2(n787), 
        .ZN(n61) );
  ND4D0 U230 ( .A1(n64), .A2(n63), .A3(n62), .A4(n61), .ZN(n65) );
  NR3D0 U231 ( .A1(n67), .A2(n66), .A3(n65), .ZN(n68) );
  ND4D0 U232 ( .A1(n71), .A2(n70), .A3(n69), .A4(n68), .ZN(B[0]) );
  CKND2D0 U233 ( .A1(n72), .A2(n73), .ZN(n226) );
  NR2D0 U234 ( .A1(dira[3]), .A2(dira[4]), .ZN(n224) );
  CKND2D0 U235 ( .A1(n224), .A2(n240), .ZN(n74) );
  NR2D0 U236 ( .A1(n226), .A2(n74), .ZN(n1121) );
  CKND2D0 U237 ( .A1(dira[1]), .A2(n72), .ZN(n232) );
  NR2D0 U238 ( .A1(n74), .A2(n232), .ZN(n1120) );
  AOI22D0 U239 ( .A1(\mem[0][20] ), .A2(n1121), .B1(\mem[2][20] ), .B2(n1120), 
        .ZN(n79) );
  CKND2D0 U240 ( .A1(dira[0]), .A2(n73), .ZN(n225) );
  NR2D0 U241 ( .A1(n74), .A2(n225), .ZN(n1123) );
  CKND2D0 U242 ( .A1(dira[0]), .A2(dira[1]), .ZN(n230) );
  NR2D0 U243 ( .A1(n74), .A2(n230), .ZN(n1122) );
  AOI22D0 U244 ( .A1(\mem[1][20] ), .A2(n1123), .B1(\mem[3][20] ), .B2(n1122), 
        .ZN(n78) );
  INVD0 U245 ( .I(dira[3]), .ZN(n88) );
  NR2D0 U246 ( .A1(dira[4]), .A2(n88), .ZN(n229) );
  CKND2D0 U247 ( .A1(n229), .A2(n240), .ZN(n75) );
  NR2D0 U248 ( .A1(n226), .A2(n75), .ZN(n1125) );
  NR2D0 U249 ( .A1(n232), .A2(n75), .ZN(n1124) );
  AOI22D0 U250 ( .A1(\mem[8][20] ), .A2(n1125), .B1(\mem[10][20] ), .B2(n1124), 
        .ZN(n77) );
  NR2D0 U251 ( .A1(n230), .A2(n75), .ZN(n1127) );
  NR2D0 U252 ( .A1(n225), .A2(n75), .ZN(n1126) );
  AOI22D0 U253 ( .A1(\mem[11][20] ), .A2(n1127), .B1(\mem[9][20] ), .B2(n1126), 
        .ZN(n76) );
  ND4D0 U254 ( .A1(n79), .A2(n78), .A3(n77), .A4(n76), .ZN(n103) );
  NR2D0 U255 ( .A1(n226), .A2(n80), .ZN(n1133) );
  NR2D0 U256 ( .A1(n232), .A2(n80), .ZN(n1132) );
  AOI22D0 U257 ( .A1(\mem[4][20] ), .A2(n1133), .B1(\mem[6][20] ), .B2(n1132), 
        .ZN(n85) );
  NR2D0 U258 ( .A1(n225), .A2(n80), .ZN(n1135) );
  NR2D0 U259 ( .A1(n230), .A2(n80), .ZN(n1134) );
  CKND2D0 U260 ( .A1(dira[2]), .A2(n229), .ZN(n81) );
  NR2D0 U261 ( .A1(n226), .A2(n81), .ZN(n1137) );
  NR2D0 U262 ( .A1(n232), .A2(n81), .ZN(n1136) );
  AOI22D0 U263 ( .A1(\mem[12][20] ), .A2(n1137), .B1(\mem[14][20] ), .B2(n1136), .ZN(n83) );
  NR2D0 U264 ( .A1(n225), .A2(n81), .ZN(n1139) );
  NR2D0 U265 ( .A1(n230), .A2(n81), .ZN(n1138) );
  AOI22D0 U266 ( .A1(\mem[13][20] ), .A2(n1139), .B1(\mem[15][20] ), .B2(n1138), .ZN(n82) );
  ND4D0 U267 ( .A1(n85), .A2(n84), .A3(n83), .A4(n82), .ZN(n102) );
  NR2D0 U268 ( .A1(dira[3]), .A2(n87), .ZN(n249) );
  CKND2D0 U269 ( .A1(n249), .A2(n240), .ZN(n86) );
  NR2D0 U270 ( .A1(n226), .A2(n86), .ZN(n1145) );
  NR2D0 U271 ( .A1(n232), .A2(n86), .ZN(n1144) );
  AOI22D0 U272 ( .A1(\mem[16][20] ), .A2(n1145), .B1(\mem[18][20] ), .B2(n1144), .ZN(n93) );
  NR2D0 U273 ( .A1(n225), .A2(n86), .ZN(n1147) );
  NR2D0 U274 ( .A1(n230), .A2(n86), .ZN(n1146) );
  AOI22D0 U275 ( .A1(\mem[17][20] ), .A2(n1147), .B1(\mem[19][20] ), .B2(n1146), .ZN(n92) );
  NR2D0 U276 ( .A1(n88), .A2(n87), .ZN(n244) );
  CKND2D0 U277 ( .A1(n244), .A2(n240), .ZN(n89) );
  NR2D0 U278 ( .A1(n226), .A2(n89), .ZN(n1149) );
  NR2D0 U279 ( .A1(n232), .A2(n89), .ZN(n1148) );
  AOI22D0 U280 ( .A1(\mem[24][20] ), .A2(n1149), .B1(\mem[26][20] ), .B2(n1148), .ZN(n91) );
  NR2D0 U281 ( .A1(n225), .A2(n89), .ZN(n1151) );
  NR2D0 U282 ( .A1(n230), .A2(n89), .ZN(n1150) );
  AOI22D0 U283 ( .A1(\mem[25][20] ), .A2(n1151), .B1(\mem[27][20] ), .B2(n1150), .ZN(n90) );
  ND4D0 U284 ( .A1(n93), .A2(n92), .A3(n91), .A4(n90), .ZN(n101) );
  CKND2D0 U285 ( .A1(dira[2]), .A2(n249), .ZN(n94) );
  NR2D0 U286 ( .A1(n226), .A2(n94), .ZN(n1157) );
  NR2D0 U287 ( .A1(n232), .A2(n94), .ZN(n1156) );
  AOI22D0 U288 ( .A1(\mem[20][20] ), .A2(n1157), .B1(\mem[22][20] ), .B2(n1156), .ZN(n99) );
  NR2D0 U289 ( .A1(n225), .A2(n94), .ZN(n1159) );
  NR2D0 U290 ( .A1(n230), .A2(n94), .ZN(n1158) );
  AOI22D0 U291 ( .A1(\mem[21][20] ), .A2(n1159), .B1(\mem[23][20] ), .B2(n1158), .ZN(n98) );
  CKND2D0 U292 ( .A1(dira[2]), .A2(n244), .ZN(n95) );
  NR2D0 U293 ( .A1(n226), .A2(n95), .ZN(n1161) );
  NR2D0 U294 ( .A1(n232), .A2(n95), .ZN(n1160) );
  AOI22D0 U295 ( .A1(\mem[28][20] ), .A2(n1161), .B1(\mem[30][20] ), .B2(n1160), .ZN(n97) );
  NR2D0 U296 ( .A1(n225), .A2(n95), .ZN(n1163) );
  NR2D0 U297 ( .A1(n230), .A2(n95), .ZN(n1162) );
  AOI22D0 U298 ( .A1(\mem[29][20] ), .A2(n1163), .B1(\mem[31][20] ), .B2(n1162), .ZN(n96) );
  ND4D0 U299 ( .A1(n99), .A2(n98), .A3(n97), .A4(n96), .ZN(n100) );
  OR4D0 U300 ( .A1(n103), .A2(n102), .A3(n101), .A4(n100), .Z(A[20]) );
  AOI22D0 U301 ( .A1(\mem[0][14] ), .A2(n1121), .B1(\mem[2][14] ), .B2(n1120), 
        .ZN(n107) );
  AOI22D0 U302 ( .A1(\mem[1][14] ), .A2(n1123), .B1(\mem[3][14] ), .B2(n1122), 
        .ZN(n106) );
  AOI22D0 U303 ( .A1(\mem[8][14] ), .A2(n1125), .B1(\mem[10][14] ), .B2(n1124), 
        .ZN(n105) );
  AOI22D0 U304 ( .A1(\mem[11][14] ), .A2(n1127), .B1(\mem[9][14] ), .B2(n1126), 
        .ZN(n104) );
  ND4D0 U305 ( .A1(n107), .A2(n106), .A3(n105), .A4(n104), .ZN(n123) );
  AOI22D0 U306 ( .A1(\mem[4][14] ), .A2(n1133), .B1(\mem[6][14] ), .B2(n1132), 
        .ZN(n111) );
  AOI22D0 U307 ( .A1(\mem[5][14] ), .A2(n1135), .B1(\mem[7][14] ), .B2(n1134), 
        .ZN(n110) );
  AOI22D0 U308 ( .A1(\mem[12][14] ), .A2(n1137), .B1(\mem[14][14] ), .B2(n1136), .ZN(n109) );
  AOI22D0 U309 ( .A1(\mem[13][14] ), .A2(n1139), .B1(\mem[15][14] ), .B2(n1138), .ZN(n108) );
  ND4D0 U310 ( .A1(n111), .A2(n110), .A3(n109), .A4(n108), .ZN(n122) );
  AOI22D0 U311 ( .A1(\mem[16][14] ), .A2(n1145), .B1(\mem[18][14] ), .B2(n1144), .ZN(n115) );
  AOI22D0 U312 ( .A1(\mem[17][14] ), .A2(n1147), .B1(\mem[19][14] ), .B2(n1146), .ZN(n114) );
  AOI22D0 U313 ( .A1(\mem[24][14] ), .A2(n1149), .B1(\mem[26][14] ), .B2(n1148), .ZN(n113) );
  AOI22D0 U314 ( .A1(\mem[25][14] ), .A2(n1151), .B1(\mem[27][14] ), .B2(n1150), .ZN(n112) );
  ND4D0 U315 ( .A1(n115), .A2(n114), .A3(n113), .A4(n112), .ZN(n121) );
  AOI22D0 U316 ( .A1(\mem[20][14] ), .A2(n1157), .B1(\mem[22][14] ), .B2(n1156), .ZN(n119) );
  AOI22D0 U317 ( .A1(\mem[21][14] ), .A2(n1159), .B1(\mem[23][14] ), .B2(n1158), .ZN(n118) );
  AOI22D0 U318 ( .A1(\mem[29][14] ), .A2(n1163), .B1(\mem[31][14] ), .B2(n1162), .ZN(n116) );
  ND4D0 U319 ( .A1(n119), .A2(n118), .A3(n117), .A4(n116), .ZN(n120) );
  OR4D0 U320 ( .A1(n123), .A2(n122), .A3(n121), .A4(n120), .Z(A[14]) );
  AOI22D0 U321 ( .A1(\mem[0][8] ), .A2(n1121), .B1(\mem[2][8] ), .B2(n1120), 
        .ZN(n127) );
  AOI22D0 U322 ( .A1(\mem[1][8] ), .A2(n1123), .B1(\mem[3][8] ), .B2(n1122), 
        .ZN(n126) );
  AOI22D0 U323 ( .A1(\mem[8][8] ), .A2(n1125), .B1(\mem[10][8] ), .B2(n1124), 
        .ZN(n125) );
  AOI22D0 U324 ( .A1(\mem[11][8] ), .A2(n1127), .B1(\mem[9][8] ), .B2(n1126), 
        .ZN(n124) );
  ND4D0 U325 ( .A1(n127), .A2(n126), .A3(n125), .A4(n124), .ZN(n143) );
  AOI22D0 U326 ( .A1(\mem[4][8] ), .A2(n1133), .B1(\mem[6][8] ), .B2(n1132), 
        .ZN(n131) );
  AOI22D0 U327 ( .A1(\mem[5][8] ), .A2(n1135), .B1(\mem[7][8] ), .B2(n1134), 
        .ZN(n130) );
  AOI22D0 U328 ( .A1(\mem[12][8] ), .A2(n1137), .B1(\mem[14][8] ), .B2(n1136), 
        .ZN(n129) );
  AOI22D0 U329 ( .A1(\mem[13][8] ), .A2(n1139), .B1(\mem[15][8] ), .B2(n1138), 
        .ZN(n128) );
  AOI22D0 U330 ( .A1(\mem[17][8] ), .A2(n1147), .B1(\mem[19][8] ), .B2(n1146), 
        .ZN(n134) );
  AOI22D0 U331 ( .A1(\mem[24][8] ), .A2(n1149), .B1(\mem[26][8] ), .B2(n1148), 
        .ZN(n133) );
  AOI22D0 U332 ( .A1(\mem[25][8] ), .A2(n1151), .B1(\mem[27][8] ), .B2(n1150), 
        .ZN(n132) );
  ND4D0 U333 ( .A1(n135), .A2(n134), .A3(n133), .A4(n132), .ZN(n141) );
  AOI22D0 U334 ( .A1(\mem[20][8] ), .A2(n1157), .B1(\mem[22][8] ), .B2(n1156), 
        .ZN(n139) );
  AOI22D0 U335 ( .A1(\mem[21][8] ), .A2(n1159), .B1(\mem[23][8] ), .B2(n1158), 
        .ZN(n138) );
  AOI22D0 U336 ( .A1(\mem[28][8] ), .A2(n1161), .B1(\mem[30][8] ), .B2(n1160), 
        .ZN(n137) );
  AOI22D0 U337 ( .A1(\mem[29][8] ), .A2(n1163), .B1(\mem[31][8] ), .B2(n1162), 
        .ZN(n136) );
  ND4D0 U338 ( .A1(n139), .A2(n138), .A3(n137), .A4(n136), .ZN(n140) );
  OR4D0 U339 ( .A1(n143), .A2(n142), .A3(n141), .A4(n140), .Z(A[8]) );
  AOI22D0 U340 ( .A1(\mem[0][5] ), .A2(n1121), .B1(\mem[2][5] ), .B2(n1120), 
        .ZN(n147) );
  AOI22D0 U341 ( .A1(\mem[1][5] ), .A2(n1123), .B1(\mem[3][5] ), .B2(n1122), 
        .ZN(n146) );
  AOI22D0 U342 ( .A1(\mem[8][5] ), .A2(n1125), .B1(\mem[10][5] ), .B2(n1124), 
        .ZN(n145) );
  AOI22D0 U343 ( .A1(\mem[11][5] ), .A2(n1127), .B1(\mem[9][5] ), .B2(n1126), 
        .ZN(n144) );
  ND4D0 U344 ( .A1(n147), .A2(n146), .A3(n145), .A4(n144), .ZN(n163) );
  AOI22D0 U345 ( .A1(\mem[4][5] ), .A2(n1133), .B1(\mem[6][5] ), .B2(n1132), 
        .ZN(n151) );
  AOI22D0 U346 ( .A1(\mem[12][5] ), .A2(n1137), .B1(\mem[14][5] ), .B2(n1136), 
        .ZN(n149) );
  AOI22D0 U347 ( .A1(\mem[13][5] ), .A2(n1139), .B1(\mem[15][5] ), .B2(n1138), 
        .ZN(n148) );
  ND4D0 U348 ( .A1(n151), .A2(n150), .A3(n149), .A4(n148), .ZN(n162) );
  AOI22D0 U349 ( .A1(\mem[16][5] ), .A2(n1145), .B1(\mem[18][5] ), .B2(n1144), 
        .ZN(n155) );
  AOI22D0 U350 ( .A1(\mem[17][5] ), .A2(n1147), .B1(\mem[19][5] ), .B2(n1146), 
        .ZN(n154) );
  AOI22D0 U351 ( .A1(\mem[24][5] ), .A2(n1149), .B1(\mem[26][5] ), .B2(n1148), 
        .ZN(n153) );
  AOI22D0 U352 ( .A1(\mem[25][5] ), .A2(n1151), .B1(\mem[27][5] ), .B2(n1150), 
        .ZN(n152) );
  ND4D0 U353 ( .A1(n155), .A2(n154), .A3(n153), .A4(n152), .ZN(n161) );
  AOI22D0 U354 ( .A1(\mem[20][5] ), .A2(n1157), .B1(\mem[22][5] ), .B2(n1156), 
        .ZN(n159) );
  AOI22D0 U355 ( .A1(\mem[21][5] ), .A2(n1159), .B1(\mem[23][5] ), .B2(n1158), 
        .ZN(n158) );
  AOI22D0 U356 ( .A1(\mem[28][5] ), .A2(n1161), .B1(\mem[30][5] ), .B2(n1160), 
        .ZN(n157) );
  AOI22D0 U357 ( .A1(\mem[29][5] ), .A2(n1163), .B1(\mem[31][5] ), .B2(n1162), 
        .ZN(n156) );
  ND4D0 U358 ( .A1(n159), .A2(n158), .A3(n157), .A4(n156), .ZN(n160) );
  OR4D0 U359 ( .A1(n163), .A2(n162), .A3(n161), .A4(n160), .Z(A[5]) );
  AOI22D0 U360 ( .A1(\mem[0][2] ), .A2(n1121), .B1(\mem[2][2] ), .B2(n1120), 
        .ZN(n167) );
  AOI22D0 U361 ( .A1(\mem[1][2] ), .A2(n1123), .B1(\mem[3][2] ), .B2(n1122), 
        .ZN(n166) );
  AOI22D0 U362 ( .A1(\mem[11][2] ), .A2(n1127), .B1(\mem[9][2] ), .B2(n1126), 
        .ZN(n164) );
  ND4D0 U363 ( .A1(n167), .A2(n166), .A3(n165), .A4(n164), .ZN(n183) );
  AOI22D0 U364 ( .A1(\mem[4][2] ), .A2(n1133), .B1(\mem[6][2] ), .B2(n1132), 
        .ZN(n171) );
  AOI22D0 U365 ( .A1(\mem[5][2] ), .A2(n1135), .B1(\mem[7][2] ), .B2(n1134), 
        .ZN(n170) );
  AOI22D0 U366 ( .A1(\mem[12][2] ), .A2(n1137), .B1(\mem[14][2] ), .B2(n1136), 
        .ZN(n169) );
  AOI22D0 U367 ( .A1(\mem[13][2] ), .A2(n1139), .B1(\mem[15][2] ), .B2(n1138), 
        .ZN(n168) );
  ND4D0 U368 ( .A1(n171), .A2(n170), .A3(n169), .A4(n168), .ZN(n182) );
  AOI22D0 U369 ( .A1(\mem[16][2] ), .A2(n1145), .B1(\mem[18][2] ), .B2(n1144), 
        .ZN(n175) );
  AOI22D0 U370 ( .A1(\mem[17][2] ), .A2(n1147), .B1(\mem[19][2] ), .B2(n1146), 
        .ZN(n174) );
  AOI22D0 U371 ( .A1(\mem[24][2] ), .A2(n1149), .B1(\mem[26][2] ), .B2(n1148), 
        .ZN(n173) );
  AOI22D0 U372 ( .A1(\mem[25][2] ), .A2(n1151), .B1(\mem[27][2] ), .B2(n1150), 
        .ZN(n172) );
  ND4D0 U373 ( .A1(n175), .A2(n174), .A3(n173), .A4(n172), .ZN(n181) );
  AOI22D0 U374 ( .A1(\mem[20][2] ), .A2(n1157), .B1(\mem[22][2] ), .B2(n1156), 
        .ZN(n179) );
  AOI22D0 U375 ( .A1(\mem[21][2] ), .A2(n1159), .B1(\mem[23][2] ), .B2(n1158), 
        .ZN(n178) );
  AOI22D0 U376 ( .A1(\mem[28][2] ), .A2(n1161), .B1(\mem[30][2] ), .B2(n1160), 
        .ZN(n177) );
  AOI22D0 U377 ( .A1(\mem[29][2] ), .A2(n1163), .B1(\mem[31][2] ), .B2(n1162), 
        .ZN(n176) );
  ND4D0 U378 ( .A1(n179), .A2(n178), .A3(n177), .A4(n176), .ZN(n180) );
  OR4D0 U379 ( .A1(n183), .A2(n182), .A3(n181), .A4(n180), .Z(A[2]) );
  AOI22D0 U380 ( .A1(\mem[0][11] ), .A2(n1121), .B1(\mem[2][11] ), .B2(n1120), 
        .ZN(n187) );
  AOI22D0 U381 ( .A1(\mem[1][11] ), .A2(n1123), .B1(\mem[3][11] ), .B2(n1122), 
        .ZN(n186) );
  AOI22D0 U382 ( .A1(\mem[8][11] ), .A2(n1125), .B1(\mem[10][11] ), .B2(n1124), 
        .ZN(n185) );
  AOI22D0 U383 ( .A1(\mem[11][11] ), .A2(n1127), .B1(\mem[9][11] ), .B2(n1126), 
        .ZN(n184) );
  ND4D0 U384 ( .A1(n187), .A2(n186), .A3(n185), .A4(n184), .ZN(n203) );
  AOI22D0 U385 ( .A1(\mem[4][11] ), .A2(n1133), .B1(\mem[6][11] ), .B2(n1132), 
        .ZN(n191) );
  AOI22D0 U386 ( .A1(\mem[5][11] ), .A2(n1135), .B1(\mem[7][11] ), .B2(n1134), 
        .ZN(n190) );
  AOI22D0 U387 ( .A1(\mem[12][11] ), .A2(n1137), .B1(\mem[14][11] ), .B2(n1136), .ZN(n189) );
  AOI22D0 U388 ( .A1(\mem[13][11] ), .A2(n1139), .B1(\mem[15][11] ), .B2(n1138), .ZN(n188) );
  ND4D0 U389 ( .A1(n191), .A2(n190), .A3(n189), .A4(n188), .ZN(n202) );
  AOI22D0 U390 ( .A1(\mem[16][11] ), .A2(n1145), .B1(\mem[18][11] ), .B2(n1144), .ZN(n195) );
  AOI22D0 U391 ( .A1(\mem[17][11] ), .A2(n1147), .B1(\mem[19][11] ), .B2(n1146), .ZN(n194) );
  AOI22D0 U392 ( .A1(\mem[24][11] ), .A2(n1149), .B1(\mem[26][11] ), .B2(n1148), .ZN(n193) );
  ND4D0 U393 ( .A1(n195), .A2(n194), .A3(n193), .A4(n192), .ZN(n201) );
  AOI22D0 U394 ( .A1(\mem[20][11] ), .A2(n1157), .B1(\mem[22][11] ), .B2(n1156), .ZN(n199) );
  AOI22D0 U395 ( .A1(\mem[21][11] ), .A2(n1159), .B1(\mem[23][11] ), .B2(n1158), .ZN(n198) );
  AOI22D0 U396 ( .A1(\mem[28][11] ), .A2(n1161), .B1(\mem[30][11] ), .B2(n1160), .ZN(n197) );
  AOI22D0 U397 ( .A1(\mem[29][11] ), .A2(n1163), .B1(\mem[31][11] ), .B2(n1162), .ZN(n196) );
  ND4D0 U398 ( .A1(n199), .A2(n198), .A3(n197), .A4(n196), .ZN(n200) );
  OR4D0 U399 ( .A1(n203), .A2(n202), .A3(n201), .A4(n200), .Z(A[11]) );
  AOI22D0 U400 ( .A1(\mem[0][17] ), .A2(n1121), .B1(\mem[2][17] ), .B2(n1120), 
        .ZN(n207) );
  AOI22D0 U401 ( .A1(\mem[1][17] ), .A2(n1123), .B1(\mem[3][17] ), .B2(n1122), 
        .ZN(n206) );
  AOI22D0 U402 ( .A1(\mem[11][17] ), .A2(n1127), .B1(\mem[9][17] ), .B2(n1126), 
        .ZN(n204) );
  ND4D0 U403 ( .A1(n207), .A2(n206), .A3(n205), .A4(n204), .ZN(n223) );
  AOI22D0 U404 ( .A1(\mem[4][17] ), .A2(n1133), .B1(\mem[6][17] ), .B2(n1132), 
        .ZN(n211) );
  AOI22D0 U405 ( .A1(\mem[5][17] ), .A2(n1135), .B1(\mem[7][17] ), .B2(n1134), 
        .ZN(n210) );
  AOI22D0 U406 ( .A1(\mem[12][17] ), .A2(n1137), .B1(\mem[14][17] ), .B2(n1136), .ZN(n209) );
  AOI22D0 U407 ( .A1(\mem[13][17] ), .A2(n1139), .B1(\mem[15][17] ), .B2(n1138), .ZN(n208) );
  ND4D0 U408 ( .A1(n211), .A2(n210), .A3(n209), .A4(n208), .ZN(n222) );
  AOI22D0 U409 ( .A1(\mem[16][17] ), .A2(n1145), .B1(\mem[18][17] ), .B2(n1144), .ZN(n215) );
  AOI22D0 U410 ( .A1(\mem[17][17] ), .A2(n1147), .B1(\mem[19][17] ), .B2(n1146), .ZN(n214) );
  AOI22D0 U411 ( .A1(\mem[24][17] ), .A2(n1149), .B1(\mem[26][17] ), .B2(n1148), .ZN(n213) );
  AOI22D0 U412 ( .A1(\mem[25][17] ), .A2(n1151), .B1(\mem[27][17] ), .B2(n1150), .ZN(n212) );
  ND4D0 U413 ( .A1(n215), .A2(n214), .A3(n213), .A4(n212), .ZN(n221) );
  AOI22D0 U414 ( .A1(\mem[20][17] ), .A2(n1157), .B1(\mem[22][17] ), .B2(n1156), .ZN(n219) );
  AOI22D0 U415 ( .A1(\mem[21][17] ), .A2(n1159), .B1(\mem[23][17] ), .B2(n1158), .ZN(n218) );
  AOI22D0 U416 ( .A1(\mem[28][17] ), .A2(n1161), .B1(\mem[30][17] ), .B2(n1160), .ZN(n217) );
  AOI22D0 U417 ( .A1(\mem[29][17] ), .A2(n1163), .B1(\mem[31][17] ), .B2(n1162), .ZN(n216) );
  ND4D0 U418 ( .A1(n219), .A2(n218), .A3(n217), .A4(n216), .ZN(n220) );
  OR4D0 U419 ( .A1(n223), .A2(n222), .A3(n221), .A4(n220), .Z(A[17]) );
  CKND2D0 U420 ( .A1(write), .A2(n224), .ZN(n242) );
  INVD0 U421 ( .I(n225), .ZN(n234) );
  CKND2D0 U422 ( .A1(n234), .A2(n240), .ZN(n275) );
  NR2XD0 U423 ( .A1(n242), .A2(n275), .ZN(n228) );
  INVD0 U424 ( .I(data[1]), .ZN(n505) );
  MAOI22D0 U425 ( .A1(n228), .A2(n505), .B1(\mem[1][1] ), .B2(n228), .ZN(n1891) );
  INVD0 U426 ( .I(data[2]), .ZN(n755) );
  MAOI22D0 U427 ( .A1(n228), .A2(n755), .B1(\mem[1][2] ), .B2(n228), .ZN(n1892) );
  INVD0 U428 ( .I(data[3]), .ZN(n483) );
  MAOI22D0 U429 ( .A1(n228), .A2(n483), .B1(\mem[1][3] ), .B2(n228), .ZN(n1893) );
  INVD0 U430 ( .I(data[4]), .ZN(n527) );
  MAOI22D0 U431 ( .A1(n228), .A2(n527), .B1(\mem[1][4] ), .B2(n228), .ZN(n1894) );
  INVD0 U432 ( .I(data[5]), .ZN(n461) );
  MAOI22D0 U433 ( .A1(n228), .A2(n461), .B1(\mem[1][5] ), .B2(n228), .ZN(n1895) );
  INVD0 U434 ( .I(data[6]), .ZN(n549) );
  MAOI22D0 U435 ( .A1(n228), .A2(n549), .B1(\mem[1][6] ), .B2(n228), .ZN(n1896) );
  INVD0 U436 ( .I(data[7]), .ZN(n439) );
  MAOI22D0 U437 ( .A1(n228), .A2(n439), .B1(\mem[1][7] ), .B2(n228), .ZN(n1897) );
  MAOI22D0 U438 ( .A1(n228), .A2(n571), .B1(\mem[1][8] ), .B2(n228), .ZN(n1898) );
  INVD0 U439 ( .I(data[9]), .ZN(n417) );
  MAOI22D0 U440 ( .A1(n228), .A2(n417), .B1(\mem[1][9] ), .B2(n228), .ZN(n1899) );
  INVD0 U441 ( .I(data[10]), .ZN(n593) );
  MAOI22D0 U442 ( .A1(n228), .A2(n593), .B1(\mem[1][10] ), .B2(n228), .ZN(
        n1900) );
  INVD0 U443 ( .I(data[11]), .ZN(n395) );
  MAOI22D0 U444 ( .A1(n228), .A2(n395), .B1(\mem[1][11] ), .B2(n228), .ZN(
        n1901) );
  INVD0 U445 ( .I(data[12]), .ZN(n615) );
  MAOI22D0 U446 ( .A1(n228), .A2(n615), .B1(\mem[1][12] ), .B2(n228), .ZN(
        n1902) );
  INVD0 U447 ( .I(data[13]), .ZN(n373) );
  MAOI22D0 U448 ( .A1(n228), .A2(n373), .B1(\mem[1][13] ), .B2(n228), .ZN(
        n1903) );
  INVD0 U449 ( .I(data[14]), .ZN(n637) );
  INVD0 U450 ( .I(data[15]), .ZN(n351) );
  MAOI22D0 U451 ( .A1(n228), .A2(n351), .B1(\mem[1][15] ), .B2(n228), .ZN(
        n1905) );
  INVD0 U452 ( .I(data[16]), .ZN(n659) );
  MAOI22D0 U453 ( .A1(n228), .A2(n659), .B1(\mem[1][16] ), .B2(n228), .ZN(
        n1906) );
  INVD0 U454 ( .I(data[17]), .ZN(n329) );
  MAOI22D0 U455 ( .A1(n228), .A2(n329), .B1(\mem[1][17] ), .B2(n228), .ZN(
        n1907) );
  INVD0 U456 ( .I(data[18]), .ZN(n681) );
  MAOI22D0 U457 ( .A1(n228), .A2(n681), .B1(\mem[1][18] ), .B2(n228), .ZN(
        n1908) );
  INVD0 U458 ( .I(data[19]), .ZN(n307) );
  MAOI22D0 U459 ( .A1(n228), .A2(n307), .B1(\mem[1][19] ), .B2(n228), .ZN(
        n1909) );
  INVD0 U460 ( .I(data[20]), .ZN(n703) );
  MAOI22D0 U461 ( .A1(n228), .A2(n703), .B1(\mem[1][20] ), .B2(n228), .ZN(
        n1910) );
  INVD0 U462 ( .I(data[21]), .ZN(n285) );
  MAOI22D0 U463 ( .A1(n228), .A2(n285), .B1(\mem[1][21] ), .B2(n228), .ZN(
        n1911) );
  INVD0 U464 ( .I(data[22]), .ZN(n725) );
  MAOI22D0 U465 ( .A1(n228), .A2(n725), .B1(\mem[1][22] ), .B2(n228), .ZN(
        n1912) );
  MAOI22D0 U466 ( .A1(n228), .A2(n279), .B1(\mem[1][23] ), .B2(n228), .ZN(
        n1913) );
  INVD0 U467 ( .I(n226), .ZN(n236) );
  CKND2D0 U468 ( .A1(n236), .A2(n240), .ZN(n278) );
  NR2XD0 U469 ( .A1(n278), .A2(n242), .ZN(n227) );
  MAOI22D0 U470 ( .A1(n227), .A2(n281), .B1(\mem[0][0] ), .B2(n227), .ZN(n1914) );
  MAOI22D0 U471 ( .A1(n227), .A2(n505), .B1(\mem[0][1] ), .B2(n227), .ZN(n1915) );
  MAOI22D0 U472 ( .A1(n227), .A2(n755), .B1(\mem[0][2] ), .B2(n227), .ZN(n1916) );
  MAOI22D0 U473 ( .A1(n227), .A2(n483), .B1(\mem[0][3] ), .B2(n227), .ZN(n1917) );
  MAOI22D0 U474 ( .A1(n227), .A2(n527), .B1(\mem[0][4] ), .B2(n227), .ZN(n1918) );
  MAOI22D0 U475 ( .A1(n227), .A2(n549), .B1(\mem[0][6] ), .B2(n227), .ZN(n1920) );
  MAOI22D0 U476 ( .A1(n227), .A2(n439), .B1(\mem[0][7] ), .B2(n227), .ZN(n1921) );
  MAOI22D0 U477 ( .A1(n227), .A2(n571), .B1(\mem[0][8] ), .B2(n227), .ZN(n1922) );
  MAOI22D0 U478 ( .A1(n227), .A2(n417), .B1(\mem[0][9] ), .B2(n227), .ZN(n1923) );
  MAOI22D0 U479 ( .A1(n227), .A2(n593), .B1(\mem[0][10] ), .B2(n227), .ZN(
        n1924) );
  MAOI22D0 U480 ( .A1(n227), .A2(n395), .B1(\mem[0][11] ), .B2(n227), .ZN(
        n1925) );
  MAOI22D0 U481 ( .A1(n227), .A2(n615), .B1(\mem[0][12] ), .B2(n227), .ZN(
        n1926) );
  MAOI22D0 U482 ( .A1(n227), .A2(n373), .B1(\mem[0][13] ), .B2(n227), .ZN(
        n1927) );
  MAOI22D0 U483 ( .A1(n227), .A2(n637), .B1(\mem[0][14] ), .B2(n227), .ZN(
        n1928) );
  MAOI22D0 U484 ( .A1(n227), .A2(n351), .B1(\mem[0][15] ), .B2(n227), .ZN(
        n1929) );
  MAOI22D0 U485 ( .A1(n227), .A2(n659), .B1(\mem[0][16] ), .B2(n227), .ZN(
        n1930) );
  MAOI22D0 U486 ( .A1(n227), .A2(n329), .B1(\mem[0][17] ), .B2(n227), .ZN(
        n1931) );
  MAOI22D0 U487 ( .A1(n227), .A2(n681), .B1(\mem[0][18] ), .B2(n227), .ZN(
        n1932) );
  MAOI22D0 U488 ( .A1(n227), .A2(n307), .B1(\mem[0][19] ), .B2(n227), .ZN(
        n1933) );
  MAOI22D0 U489 ( .A1(n227), .A2(n285), .B1(\mem[0][21] ), .B2(n227), .ZN(
        n1935) );
  MAOI22D0 U490 ( .A1(n227), .A2(n725), .B1(\mem[0][22] ), .B2(n227), .ZN(
        n1936) );
  MAOI22D0 U491 ( .A1(n227), .A2(n279), .B1(\mem[0][23] ), .B2(n227), .ZN(
        n1937) );
  MAOI22D0 U492 ( .A1(n228), .A2(n281), .B1(\mem[1][0] ), .B2(n228), .ZN(n1890) );
  CKND2D0 U493 ( .A1(write), .A2(n229), .ZN(n265) );
  NR2XD0 U494 ( .A1(n278), .A2(n265), .ZN(n267) );
  MAOI22D0 U495 ( .A1(n267), .A2(n615), .B1(\mem[8][12] ), .B2(n267), .ZN(
        n1734) );
  MAOI22D0 U496 ( .A1(n267), .A2(n373), .B1(\mem[8][13] ), .B2(n267), .ZN(
        n1735) );
  MAOI22D0 U497 ( .A1(n267), .A2(n637), .B1(\mem[8][14] ), .B2(n267), .ZN(
        n1736) );
  MAOI22D0 U498 ( .A1(n267), .A2(n351), .B1(\mem[8][15] ), .B2(n267), .ZN(
        n1737) );
  MAOI22D0 U499 ( .A1(n267), .A2(n659), .B1(\mem[8][16] ), .B2(n267), .ZN(
        n1738) );
  MAOI22D0 U500 ( .A1(n267), .A2(n681), .B1(\mem[8][18] ), .B2(n267), .ZN(
        n1740) );
  MAOI22D0 U501 ( .A1(n267), .A2(n307), .B1(\mem[8][19] ), .B2(n267), .ZN(
        n1741) );
  MAOI22D0 U502 ( .A1(n267), .A2(n703), .B1(\mem[8][20] ), .B2(n267), .ZN(
        n1742) );
  MAOI22D0 U503 ( .A1(n267), .A2(n285), .B1(\mem[8][21] ), .B2(n267), .ZN(
        n1743) );
  MAOI22D0 U504 ( .A1(n267), .A2(n725), .B1(\mem[8][22] ), .B2(n267), .ZN(
        n1744) );
  MAOI22D0 U505 ( .A1(n267), .A2(n279), .B1(\mem[8][23] ), .B2(n267), .ZN(
        n1745) );
  INVD0 U506 ( .I(n230), .ZN(n238) );
  CKND2D0 U507 ( .A1(dira[2]), .A2(n238), .ZN(n257) );
  NR2XD0 U508 ( .A1(n242), .A2(n257), .ZN(n231) );
  MAOI22D0 U509 ( .A1(n231), .A2(n281), .B1(\mem[7][0] ), .B2(n231), .ZN(n1746) );
  MAOI22D0 U510 ( .A1(n231), .A2(n505), .B1(\mem[7][1] ), .B2(n231), .ZN(n1747) );
  MAOI22D0 U511 ( .A1(n231), .A2(n755), .B1(\mem[7][2] ), .B2(n231), .ZN(n1748) );
  MAOI22D0 U512 ( .A1(n231), .A2(n483), .B1(\mem[7][3] ), .B2(n231), .ZN(n1749) );
  MAOI22D0 U513 ( .A1(n231), .A2(n527), .B1(\mem[7][4] ), .B2(n231), .ZN(n1750) );
  MAOI22D0 U514 ( .A1(n231), .A2(n461), .B1(\mem[7][5] ), .B2(n231), .ZN(n1751) );
  MAOI22D0 U515 ( .A1(n231), .A2(n549), .B1(\mem[7][6] ), .B2(n231), .ZN(n1752) );
  MAOI22D0 U516 ( .A1(n231), .A2(n439), .B1(\mem[7][7] ), .B2(n231), .ZN(n1753) );
  MAOI22D0 U517 ( .A1(n231), .A2(n417), .B1(\mem[7][9] ), .B2(n231), .ZN(n1755) );
  MAOI22D0 U518 ( .A1(n231), .A2(n593), .B1(\mem[7][10] ), .B2(n231), .ZN(
        n1756) );
  MAOI22D0 U519 ( .A1(n231), .A2(n395), .B1(\mem[7][11] ), .B2(n231), .ZN(
        n1757) );
  MAOI22D0 U520 ( .A1(n231), .A2(n615), .B1(\mem[7][12] ), .B2(n231), .ZN(
        n1758) );
  MAOI22D0 U521 ( .A1(n231), .A2(n373), .B1(\mem[7][13] ), .B2(n231), .ZN(
        n1759) );
  MAOI22D0 U522 ( .A1(n231), .A2(n637), .B1(\mem[7][14] ), .B2(n231), .ZN(
        n1760) );
  MAOI22D0 U523 ( .A1(n231), .A2(n351), .B1(\mem[7][15] ), .B2(n231), .ZN(
        n1761) );
  MAOI22D0 U524 ( .A1(n231), .A2(n659), .B1(\mem[7][16] ), .B2(n231), .ZN(
        n1762) );
  MAOI22D0 U525 ( .A1(n231), .A2(n329), .B1(\mem[7][17] ), .B2(n231), .ZN(
        n1763) );
  MAOI22D0 U526 ( .A1(n231), .A2(n681), .B1(\mem[7][18] ), .B2(n231), .ZN(
        n1764) );
  MAOI22D0 U527 ( .A1(n231), .A2(n307), .B1(\mem[7][19] ), .B2(n231), .ZN(
        n1765) );
  MAOI22D0 U528 ( .A1(n231), .A2(n703), .B1(\mem[7][20] ), .B2(n231), .ZN(
        n1766) );
  MAOI22D0 U529 ( .A1(n231), .A2(n285), .B1(\mem[7][21] ), .B2(n231), .ZN(
        n1767) );
  MAOI22D0 U530 ( .A1(n231), .A2(n725), .B1(\mem[7][22] ), .B2(n231), .ZN(
        n1768) );
  INVD0 U531 ( .I(n232), .ZN(n241) );
  CKND2D0 U532 ( .A1(dira[2]), .A2(n241), .ZN(n258) );
  NR2XD0 U533 ( .A1(n242), .A2(n258), .ZN(n233) );
  MAOI22D0 U534 ( .A1(n233), .A2(n281), .B1(\mem[6][0] ), .B2(n233), .ZN(n1770) );
  MAOI22D0 U535 ( .A1(n233), .A2(n505), .B1(\mem[6][1] ), .B2(n233), .ZN(n1771) );
  MAOI22D0 U536 ( .A1(n233), .A2(n755), .B1(\mem[6][2] ), .B2(n233), .ZN(n1772) );
  MAOI22D0 U537 ( .A1(n233), .A2(n483), .B1(\mem[6][3] ), .B2(n233), .ZN(n1773) );
  MAOI22D0 U538 ( .A1(n233), .A2(n527), .B1(\mem[6][4] ), .B2(n233), .ZN(n1774) );
  MAOI22D0 U539 ( .A1(n233), .A2(n461), .B1(\mem[6][5] ), .B2(n233), .ZN(n1775) );
  MAOI22D0 U540 ( .A1(n233), .A2(n549), .B1(\mem[6][6] ), .B2(n233), .ZN(n1776) );
  MAOI22D0 U541 ( .A1(n233), .A2(n439), .B1(\mem[6][7] ), .B2(n233), .ZN(n1777) );
  MAOI22D0 U542 ( .A1(n233), .A2(n571), .B1(\mem[6][8] ), .B2(n233), .ZN(n1778) );
  MAOI22D0 U543 ( .A1(n233), .A2(n417), .B1(\mem[6][9] ), .B2(n233), .ZN(n1779) );
  MAOI22D0 U544 ( .A1(n233), .A2(n593), .B1(\mem[6][10] ), .B2(n233), .ZN(
        n1780) );
  MAOI22D0 U545 ( .A1(n233), .A2(n395), .B1(\mem[6][11] ), .B2(n233), .ZN(
        n1781) );
  MAOI22D0 U546 ( .A1(n233), .A2(n615), .B1(\mem[6][12] ), .B2(n233), .ZN(
        n1782) );
  MAOI22D0 U547 ( .A1(n233), .A2(n373), .B1(\mem[6][13] ), .B2(n233), .ZN(
        n1783) );
  MAOI22D0 U548 ( .A1(n233), .A2(n351), .B1(\mem[6][15] ), .B2(n233), .ZN(
        n1785) );
  MAOI22D0 U549 ( .A1(n233), .A2(n659), .B1(\mem[6][16] ), .B2(n233), .ZN(
        n1786) );
  MAOI22D0 U550 ( .A1(n233), .A2(n329), .B1(\mem[6][17] ), .B2(n233), .ZN(
        n1787) );
  MAOI22D0 U551 ( .A1(n233), .A2(n681), .B1(\mem[6][18] ), .B2(n233), .ZN(
        n1788) );
  MAOI22D0 U552 ( .A1(n233), .A2(n307), .B1(\mem[6][19] ), .B2(n233), .ZN(
        n1789) );
  MAOI22D0 U553 ( .A1(n233), .A2(n703), .B1(\mem[6][20] ), .B2(n233), .ZN(
        n1790) );
  MAOI22D0 U554 ( .A1(n233), .A2(n285), .B1(\mem[6][21] ), .B2(n233), .ZN(
        n1791) );
  MAOI22D0 U555 ( .A1(n233), .A2(n725), .B1(\mem[6][22] ), .B2(n233), .ZN(
        n1792) );
  MAOI22D0 U556 ( .A1(n233), .A2(n279), .B1(\mem[6][23] ), .B2(n233), .ZN(
        n1793) );
  CKND2D0 U557 ( .A1(dira[2]), .A2(n234), .ZN(n260) );
  NR2XD0 U558 ( .A1(n242), .A2(n260), .ZN(n235) );
  MAOI22D0 U559 ( .A1(n235), .A2(n281), .B1(\mem[5][0] ), .B2(n235), .ZN(n1794) );
  MAOI22D0 U560 ( .A1(n235), .A2(n505), .B1(\mem[5][1] ), .B2(n235), .ZN(n1795) );
  MAOI22D0 U561 ( .A1(n235), .A2(n755), .B1(\mem[5][2] ), .B2(n235), .ZN(n1796) );
  MAOI22D0 U562 ( .A1(n235), .A2(n483), .B1(\mem[5][3] ), .B2(n235), .ZN(n1797) );
  MAOI22D0 U563 ( .A1(n235), .A2(n527), .B1(\mem[5][4] ), .B2(n235), .ZN(n1798) );
  MAOI22D0 U564 ( .A1(n235), .A2(n549), .B1(\mem[5][6] ), .B2(n235), .ZN(n1800) );
  MAOI22D0 U565 ( .A1(n235), .A2(n439), .B1(\mem[5][7] ), .B2(n235), .ZN(n1801) );
  MAOI22D0 U566 ( .A1(n235), .A2(n571), .B1(\mem[5][8] ), .B2(n235), .ZN(n1802) );
  MAOI22D0 U567 ( .A1(n235), .A2(n417), .B1(\mem[5][9] ), .B2(n235), .ZN(n1803) );
  MAOI22D0 U568 ( .A1(n235), .A2(n593), .B1(\mem[5][10] ), .B2(n235), .ZN(
        n1804) );
  MAOI22D0 U569 ( .A1(n235), .A2(n395), .B1(\mem[5][11] ), .B2(n235), .ZN(
        n1805) );
  MAOI22D0 U570 ( .A1(n235), .A2(n615), .B1(\mem[5][12] ), .B2(n235), .ZN(
        n1806) );
  MAOI22D0 U571 ( .A1(n235), .A2(n373), .B1(\mem[5][13] ), .B2(n235), .ZN(
        n1807) );
  MAOI22D0 U572 ( .A1(n235), .A2(n637), .B1(\mem[5][14] ), .B2(n235), .ZN(
        n1808) );
  MAOI22D0 U573 ( .A1(n235), .A2(n351), .B1(\mem[5][15] ), .B2(n235), .ZN(
        n1809) );
  MAOI22D0 U574 ( .A1(n235), .A2(n659), .B1(\mem[5][16] ), .B2(n235), .ZN(
        n1810) );
  MAOI22D0 U575 ( .A1(n235), .A2(n329), .B1(\mem[5][17] ), .B2(n235), .ZN(
        n1811) );
  MAOI22D0 U576 ( .A1(n267), .A2(n395), .B1(\mem[8][11] ), .B2(n267), .ZN(
        n1733) );
  MAOI22D0 U577 ( .A1(n235), .A2(n681), .B1(\mem[5][18] ), .B2(n235), .ZN(
        n1812) );
  MAOI22D0 U578 ( .A1(n235), .A2(n307), .B1(\mem[5][19] ), .B2(n235), .ZN(
        n1813) );
  MAOI22D0 U579 ( .A1(n235), .A2(n285), .B1(\mem[5][21] ), .B2(n235), .ZN(
        n1815) );
  MAOI22D0 U580 ( .A1(n235), .A2(n725), .B1(\mem[5][22] ), .B2(n235), .ZN(
        n1816) );
  MAOI22D0 U581 ( .A1(n235), .A2(n279), .B1(\mem[5][23] ), .B2(n235), .ZN(
        n1817) );
  CKND2D0 U582 ( .A1(dira[2]), .A2(n236), .ZN(n268) );
  NR2XD0 U583 ( .A1(n242), .A2(n268), .ZN(n237) );
  MAOI22D0 U584 ( .A1(n237), .A2(n281), .B1(\mem[4][0] ), .B2(n237), .ZN(n1818) );
  MAOI22D0 U585 ( .A1(n237), .A2(n505), .B1(\mem[4][1] ), .B2(n237), .ZN(n1819) );
  MAOI22D0 U586 ( .A1(n237), .A2(n755), .B1(\mem[4][2] ), .B2(n237), .ZN(n1820) );
  MAOI22D0 U587 ( .A1(n237), .A2(n483), .B1(\mem[4][3] ), .B2(n237), .ZN(n1821) );
  MAOI22D0 U588 ( .A1(n237), .A2(n527), .B1(\mem[4][4] ), .B2(n237), .ZN(n1822) );
  MAOI22D0 U589 ( .A1(n237), .A2(n461), .B1(\mem[4][5] ), .B2(n237), .ZN(n1823) );
  MAOI22D0 U590 ( .A1(n237), .A2(n549), .B1(\mem[4][6] ), .B2(n237), .ZN(n1824) );
  MAOI22D0 U591 ( .A1(n237), .A2(n439), .B1(\mem[4][7] ), .B2(n237), .ZN(n1825) );
  MAOI22D0 U592 ( .A1(n237), .A2(n571), .B1(\mem[4][8] ), .B2(n237), .ZN(n1826) );
  MAOI22D0 U593 ( .A1(n237), .A2(n417), .B1(\mem[4][9] ), .B2(n237), .ZN(n1827) );
  MAOI22D0 U594 ( .A1(n237), .A2(n593), .B1(\mem[4][10] ), .B2(n237), .ZN(
        n1828) );
  MAOI22D0 U595 ( .A1(n237), .A2(n615), .B1(\mem[4][12] ), .B2(n237), .ZN(
        n1830) );
  MAOI22D0 U596 ( .A1(n237), .A2(n373), .B1(\mem[4][13] ), .B2(n237), .ZN(
        n1831) );
  MAOI22D0 U597 ( .A1(n237), .A2(n637), .B1(\mem[4][14] ), .B2(n237), .ZN(
        n1832) );
  MAOI22D0 U598 ( .A1(n237), .A2(n351), .B1(\mem[4][15] ), .B2(n237), .ZN(
        n1833) );
  MAOI22D0 U599 ( .A1(n237), .A2(n659), .B1(\mem[4][16] ), .B2(n237), .ZN(
        n1834) );
  MAOI22D0 U600 ( .A1(n237), .A2(n329), .B1(\mem[4][17] ), .B2(n237), .ZN(
        n1835) );
  MAOI22D0 U601 ( .A1(n237), .A2(n681), .B1(\mem[4][18] ), .B2(n237), .ZN(
        n1836) );
  MAOI22D0 U602 ( .A1(n237), .A2(n307), .B1(\mem[4][19] ), .B2(n237), .ZN(
        n1837) );
  MAOI22D0 U603 ( .A1(n237), .A2(n703), .B1(\mem[4][20] ), .B2(n237), .ZN(
        n1838) );
  MAOI22D0 U604 ( .A1(n237), .A2(n285), .B1(\mem[4][21] ), .B2(n237), .ZN(
        n1839) );
  MAOI22D0 U605 ( .A1(n237), .A2(n725), .B1(\mem[4][22] ), .B2(n237), .ZN(
        n1840) );
  MAOI22D0 U606 ( .A1(n237), .A2(n279), .B1(\mem[4][23] ), .B2(n237), .ZN(
        n1841) );
  CKND2D0 U607 ( .A1(n238), .A2(n240), .ZN(n270) );
  NR2XD0 U608 ( .A1(n242), .A2(n270), .ZN(n239) );
  MAOI22D0 U609 ( .A1(n239), .A2(n281), .B1(\mem[3][0] ), .B2(n239), .ZN(n1842) );
  MAOI22D0 U610 ( .A1(n239), .A2(n505), .B1(\mem[3][1] ), .B2(n239), .ZN(n1843) );
  MAOI22D0 U611 ( .A1(n239), .A2(n483), .B1(\mem[3][3] ), .B2(n239), .ZN(n1845) );
  MAOI22D0 U612 ( .A1(n239), .A2(n527), .B1(\mem[3][4] ), .B2(n239), .ZN(n1846) );
  MAOI22D0 U613 ( .A1(n239), .A2(n461), .B1(\mem[3][5] ), .B2(n239), .ZN(n1847) );
  MAOI22D0 U614 ( .A1(n239), .A2(n549), .B1(\mem[3][6] ), .B2(n239), .ZN(n1848) );
  MAOI22D0 U615 ( .A1(n239), .A2(n439), .B1(\mem[3][7] ), .B2(n239), .ZN(n1849) );
  MAOI22D0 U616 ( .A1(n239), .A2(n571), .B1(\mem[3][8] ), .B2(n239), .ZN(n1850) );
  MAOI22D0 U617 ( .A1(n239), .A2(n417), .B1(\mem[3][9] ), .B2(n239), .ZN(n1851) );
  MAOI22D0 U618 ( .A1(n239), .A2(n593), .B1(\mem[3][10] ), .B2(n239), .ZN(
        n1852) );
  MAOI22D0 U619 ( .A1(n239), .A2(n395), .B1(\mem[3][11] ), .B2(n239), .ZN(
        n1853) );
  MAOI22D0 U620 ( .A1(n239), .A2(n615), .B1(\mem[3][12] ), .B2(n239), .ZN(
        n1854) );
  MAOI22D0 U621 ( .A1(n239), .A2(n373), .B1(\mem[3][13] ), .B2(n239), .ZN(
        n1855) );
  MAOI22D0 U622 ( .A1(n239), .A2(n637), .B1(\mem[3][14] ), .B2(n239), .ZN(
        n1856) );
  MAOI22D0 U623 ( .A1(n239), .A2(n351), .B1(\mem[3][15] ), .B2(n239), .ZN(
        n1857) );
  MAOI22D0 U624 ( .A1(n239), .A2(n659), .B1(\mem[3][16] ), .B2(n239), .ZN(
        n1858) );
  MAOI22D0 U625 ( .A1(n239), .A2(n681), .B1(\mem[3][18] ), .B2(n239), .ZN(
        n1860) );
  MAOI22D0 U626 ( .A1(n239), .A2(n307), .B1(\mem[3][19] ), .B2(n239), .ZN(
        n1861) );
  MAOI22D0 U627 ( .A1(n239), .A2(n703), .B1(\mem[3][20] ), .B2(n239), .ZN(
        n1862) );
  MAOI22D0 U628 ( .A1(n239), .A2(n285), .B1(\mem[3][21] ), .B2(n239), .ZN(
        n1863) );
  MAOI22D0 U629 ( .A1(n239), .A2(n725), .B1(\mem[3][22] ), .B2(n239), .ZN(
        n1864) );
  MAOI22D0 U630 ( .A1(n239), .A2(n279), .B1(\mem[3][23] ), .B2(n239), .ZN(
        n1865) );
  CKND2D0 U631 ( .A1(n241), .A2(n240), .ZN(n272) );
  NR2XD0 U632 ( .A1(n242), .A2(n272), .ZN(n243) );
  MAOI22D0 U633 ( .A1(n243), .A2(n281), .B1(\mem[2][0] ), .B2(n243), .ZN(n1866) );
  MAOI22D0 U634 ( .A1(n243), .A2(n505), .B1(\mem[2][1] ), .B2(n243), .ZN(n1867) );
  MAOI22D0 U635 ( .A1(n243), .A2(n755), .B1(\mem[2][2] ), .B2(n243), .ZN(n1868) );
  MAOI22D0 U636 ( .A1(n243), .A2(n483), .B1(\mem[2][3] ), .B2(n243), .ZN(n1869) );
  MAOI22D0 U637 ( .A1(n243), .A2(n527), .B1(\mem[2][4] ), .B2(n243), .ZN(n1870) );
  MAOI22D0 U638 ( .A1(n243), .A2(n461), .B1(\mem[2][5] ), .B2(n243), .ZN(n1871) );
  MAOI22D0 U639 ( .A1(n243), .A2(n549), .B1(\mem[2][6] ), .B2(n243), .ZN(n1872) );
  MAOI22D0 U640 ( .A1(n243), .A2(n439), .B1(\mem[2][7] ), .B2(n243), .ZN(n1873) );
  MAOI22D0 U641 ( .A1(n243), .A2(n417), .B1(\mem[2][9] ), .B2(n243), .ZN(n1875) );
  MAOI22D0 U642 ( .A1(n243), .A2(n593), .B1(\mem[2][10] ), .B2(n243), .ZN(
        n1876) );
  MAOI22D0 U643 ( .A1(n243), .A2(n395), .B1(\mem[2][11] ), .B2(n243), .ZN(
        n1877) );
  MAOI22D0 U644 ( .A1(n243), .A2(n615), .B1(\mem[2][12] ), .B2(n243), .ZN(
        n1878) );
  MAOI22D0 U645 ( .A1(n243), .A2(n373), .B1(\mem[2][13] ), .B2(n243), .ZN(
        n1879) );
  MAOI22D0 U646 ( .A1(n243), .A2(n637), .B1(\mem[2][14] ), .B2(n243), .ZN(
        n1880) );
  MAOI22D0 U647 ( .A1(n243), .A2(n351), .B1(\mem[2][15] ), .B2(n243), .ZN(
        n1881) );
  MAOI22D0 U648 ( .A1(n243), .A2(n659), .B1(\mem[2][16] ), .B2(n243), .ZN(
        n1882) );
  MAOI22D0 U649 ( .A1(n243), .A2(n329), .B1(\mem[2][17] ), .B2(n243), .ZN(
        n1883) );
  MAOI22D0 U650 ( .A1(n243), .A2(n681), .B1(\mem[2][18] ), .B2(n243), .ZN(
        n1884) );
  MAOI22D0 U651 ( .A1(n243), .A2(n307), .B1(\mem[2][19] ), .B2(n243), .ZN(
        n1885) );
  MAOI22D0 U652 ( .A1(n243), .A2(n703), .B1(\mem[2][20] ), .B2(n243), .ZN(
        n1886) );
  MAOI22D0 U653 ( .A1(n243), .A2(n285), .B1(\mem[2][21] ), .B2(n243), .ZN(
        n1887) );
  MAOI22D0 U654 ( .A1(n243), .A2(n725), .B1(\mem[2][22] ), .B2(n243), .ZN(
        n1888) );
  MAOI22D0 U655 ( .A1(n267), .A2(n593), .B1(\mem[8][10] ), .B2(n267), .ZN(
        n1732) );
  MAOI22D0 U656 ( .A1(n267), .A2(n417), .B1(\mem[8][9] ), .B2(n267), .ZN(n1731) );
  CKND2D0 U657 ( .A1(write), .A2(n244), .ZN(n254) );
  NR2XD0 U658 ( .A1(n268), .A2(n254), .ZN(n256) );
  MAOI22D0 U659 ( .A1(n256), .A2(n681), .B1(\mem[28][18] ), .B2(n256), .ZN(
        n1260) );
  MAOI22D0 U660 ( .A1(n256), .A2(n307), .B1(\mem[28][19] ), .B2(n256), .ZN(
        n1261) );
  MAOI22D0 U661 ( .A1(n256), .A2(n703), .B1(\mem[28][20] ), .B2(n256), .ZN(
        n1262) );
  MAOI22D0 U662 ( .A1(n256), .A2(n285), .B1(\mem[28][21] ), .B2(n256), .ZN(
        n1263) );
  MAOI22D0 U663 ( .A1(n256), .A2(n725), .B1(\mem[28][22] ), .B2(n256), .ZN(
        n1264) );
  MAOI22D0 U664 ( .A1(n256), .A2(n279), .B1(\mem[28][23] ), .B2(n256), .ZN(
        n1265) );
  NR2XD0 U665 ( .A1(n270), .A2(n254), .ZN(n245) );
  MAOI22D0 U666 ( .A1(n245), .A2(n281), .B1(\mem[27][0] ), .B2(n245), .ZN(
        n1266) );
  MAOI22D0 U667 ( .A1(n245), .A2(n505), .B1(\mem[27][1] ), .B2(n245), .ZN(
        n1267) );
  MAOI22D0 U668 ( .A1(n245), .A2(n755), .B1(\mem[27][2] ), .B2(n245), .ZN(
        n1268) );
  MAOI22D0 U669 ( .A1(n245), .A2(n483), .B1(\mem[27][3] ), .B2(n245), .ZN(
        n1269) );
  MAOI22D0 U670 ( .A1(n245), .A2(n527), .B1(\mem[27][4] ), .B2(n245), .ZN(
        n1270) );
  MAOI22D0 U671 ( .A1(n245), .A2(n461), .B1(\mem[27][5] ), .B2(n245), .ZN(
        n1271) );
  MAOI22D0 U672 ( .A1(n245), .A2(n549), .B1(\mem[27][6] ), .B2(n245), .ZN(
        n1272) );
  MAOI22D0 U673 ( .A1(n245), .A2(n439), .B1(\mem[27][7] ), .B2(n245), .ZN(
        n1273) );
  MAOI22D0 U674 ( .A1(n245), .A2(n417), .B1(\mem[27][9] ), .B2(n245), .ZN(
        n1275) );
  MAOI22D0 U675 ( .A1(n245), .A2(n593), .B1(\mem[27][10] ), .B2(n245), .ZN(
        n1276) );
  MAOI22D0 U676 ( .A1(n245), .A2(n395), .B1(\mem[27][11] ), .B2(n245), .ZN(
        n1277) );
  MAOI22D0 U677 ( .A1(n245), .A2(n615), .B1(\mem[27][12] ), .B2(n245), .ZN(
        n1278) );
  MAOI22D0 U678 ( .A1(n245), .A2(n373), .B1(\mem[27][13] ), .B2(n245), .ZN(
        n1279) );
  MAOI22D0 U679 ( .A1(n245), .A2(n637), .B1(\mem[27][14] ), .B2(n245), .ZN(
        n1280) );
  MAOI22D0 U680 ( .A1(n245), .A2(n351), .B1(\mem[27][15] ), .B2(n245), .ZN(
        n1281) );
  MAOI22D0 U681 ( .A1(n245), .A2(n659), .B1(\mem[27][16] ), .B2(n245), .ZN(
        n1282) );
  MAOI22D0 U682 ( .A1(n245), .A2(n329), .B1(\mem[27][17] ), .B2(n245), .ZN(
        n1283) );
  MAOI22D0 U683 ( .A1(n245), .A2(n681), .B1(\mem[27][18] ), .B2(n245), .ZN(
        n1284) );
  MAOI22D0 U684 ( .A1(n245), .A2(n307), .B1(\mem[27][19] ), .B2(n245), .ZN(
        n1285) );
  MAOI22D0 U685 ( .A1(n245), .A2(n703), .B1(\mem[27][20] ), .B2(n245), .ZN(
        n1286) );
  MAOI22D0 U686 ( .A1(n245), .A2(n285), .B1(\mem[27][21] ), .B2(n245), .ZN(
        n1287) );
  MAOI22D0 U687 ( .A1(n245), .A2(n725), .B1(\mem[27][22] ), .B2(n245), .ZN(
        n1288) );
  NR2XD0 U688 ( .A1(n272), .A2(n254), .ZN(n246) );
  MAOI22D0 U689 ( .A1(n246), .A2(n281), .B1(\mem[26][0] ), .B2(n246), .ZN(
        n1290) );
  MAOI22D0 U690 ( .A1(n246), .A2(n505), .B1(\mem[26][1] ), .B2(n246), .ZN(
        n1291) );
  MAOI22D0 U691 ( .A1(n246), .A2(n755), .B1(\mem[26][2] ), .B2(n246), .ZN(
        n1292) );
  MAOI22D0 U692 ( .A1(n246), .A2(n483), .B1(\mem[26][3] ), .B2(n246), .ZN(
        n1293) );
  MAOI22D0 U693 ( .A1(n246), .A2(n527), .B1(\mem[26][4] ), .B2(n246), .ZN(
        n1294) );
  MAOI22D0 U694 ( .A1(n246), .A2(n461), .B1(\mem[26][5] ), .B2(n246), .ZN(
        n1295) );
  MAOI22D0 U695 ( .A1(n246), .A2(n549), .B1(\mem[26][6] ), .B2(n246), .ZN(
        n1296) );
  MAOI22D0 U696 ( .A1(n246), .A2(n439), .B1(\mem[26][7] ), .B2(n246), .ZN(
        n1297) );
  MAOI22D0 U697 ( .A1(n246), .A2(n571), .B1(\mem[26][8] ), .B2(n246), .ZN(
        n1298) );
  MAOI22D0 U698 ( .A1(n246), .A2(n417), .B1(\mem[26][9] ), .B2(n246), .ZN(
        n1299) );
  MAOI22D0 U699 ( .A1(n246), .A2(n593), .B1(\mem[26][10] ), .B2(n246), .ZN(
        n1300) );
  MAOI22D0 U700 ( .A1(n246), .A2(n395), .B1(\mem[26][11] ), .B2(n246), .ZN(
        n1301) );
  MAOI22D0 U701 ( .A1(n246), .A2(n615), .B1(\mem[26][12] ), .B2(n246), .ZN(
        n1302) );
  MAOI22D0 U702 ( .A1(n246), .A2(n373), .B1(\mem[26][13] ), .B2(n246), .ZN(
        n1303) );
  MAOI22D0 U703 ( .A1(n246), .A2(n351), .B1(\mem[26][15] ), .B2(n246), .ZN(
        n1305) );
  MAOI22D0 U704 ( .A1(n246), .A2(n659), .B1(\mem[26][16] ), .B2(n246), .ZN(
        n1306) );
  MAOI22D0 U705 ( .A1(n246), .A2(n329), .B1(\mem[26][17] ), .B2(n246), .ZN(
        n1307) );
  MAOI22D0 U706 ( .A1(n246), .A2(n681), .B1(\mem[26][18] ), .B2(n246), .ZN(
        n1308) );
  MAOI22D0 U707 ( .A1(n246), .A2(n307), .B1(\mem[26][19] ), .B2(n246), .ZN(
        n1309) );
  MAOI22D0 U708 ( .A1(n246), .A2(n703), .B1(\mem[26][20] ), .B2(n246), .ZN(
        n1310) );
  MAOI22D0 U709 ( .A1(n246), .A2(n285), .B1(\mem[26][21] ), .B2(n246), .ZN(
        n1311) );
  MAOI22D0 U710 ( .A1(n246), .A2(n725), .B1(\mem[26][22] ), .B2(n246), .ZN(
        n1312) );
  MAOI22D0 U711 ( .A1(n246), .A2(n279), .B1(\mem[26][23] ), .B2(n246), .ZN(
        n1313) );
  NR2XD0 U712 ( .A1(n275), .A2(n254), .ZN(n247) );
  MAOI22D0 U713 ( .A1(n247), .A2(n281), .B1(\mem[25][0] ), .B2(n247), .ZN(
        n1314) );
  MAOI22D0 U714 ( .A1(n247), .A2(n505), .B1(\mem[25][1] ), .B2(n247), .ZN(
        n1315) );
  MAOI22D0 U715 ( .A1(n247), .A2(n755), .B1(\mem[25][2] ), .B2(n247), .ZN(
        n1316) );
  MAOI22D0 U716 ( .A1(n247), .A2(n483), .B1(\mem[25][3] ), .B2(n247), .ZN(
        n1317) );
  MAOI22D0 U717 ( .A1(n247), .A2(n527), .B1(\mem[25][4] ), .B2(n247), .ZN(
        n1318) );
  MAOI22D0 U718 ( .A1(n247), .A2(n549), .B1(\mem[25][6] ), .B2(n247), .ZN(
        n1320) );
  MAOI22D0 U719 ( .A1(n247), .A2(n439), .B1(\mem[25][7] ), .B2(n247), .ZN(
        n1321) );
  MAOI22D0 U720 ( .A1(n247), .A2(n571), .B1(\mem[25][8] ), .B2(n247), .ZN(
        n1322) );
  MAOI22D0 U721 ( .A1(n247), .A2(n417), .B1(\mem[25][9] ), .B2(n247), .ZN(
        n1323) );
  MAOI22D0 U722 ( .A1(n247), .A2(n593), .B1(\mem[25][10] ), .B2(n247), .ZN(
        n1324) );
  MAOI22D0 U723 ( .A1(n247), .A2(n395), .B1(\mem[25][11] ), .B2(n247), .ZN(
        n1325) );
  MAOI22D0 U724 ( .A1(n247), .A2(n615), .B1(\mem[25][12] ), .B2(n247), .ZN(
        n1326) );
  MAOI22D0 U725 ( .A1(n247), .A2(n373), .B1(\mem[25][13] ), .B2(n247), .ZN(
        n1327) );
  MAOI22D0 U726 ( .A1(n247), .A2(n637), .B1(\mem[25][14] ), .B2(n247), .ZN(
        n1328) );
  MAOI22D0 U727 ( .A1(n247), .A2(n351), .B1(\mem[25][15] ), .B2(n247), .ZN(
        n1329) );
  MAOI22D0 U728 ( .A1(n247), .A2(n659), .B1(\mem[25][16] ), .B2(n247), .ZN(
        n1330) );
  MAOI22D0 U729 ( .A1(n247), .A2(n329), .B1(\mem[25][17] ), .B2(n247), .ZN(
        n1331) );
  MAOI22D0 U730 ( .A1(n247), .A2(n681), .B1(\mem[25][18] ), .B2(n247), .ZN(
        n1332) );
  MAOI22D0 U731 ( .A1(n247), .A2(n307), .B1(\mem[25][19] ), .B2(n247), .ZN(
        n1333) );
  MAOI22D0 U732 ( .A1(n247), .A2(n285), .B1(\mem[25][21] ), .B2(n247), .ZN(
        n1335) );
  MAOI22D0 U733 ( .A1(n247), .A2(n725), .B1(\mem[25][22] ), .B2(n247), .ZN(
        n1336) );
  MAOI22D0 U734 ( .A1(n256), .A2(n659), .B1(\mem[28][16] ), .B2(n256), .ZN(
        n1258) );
  MAOI22D0 U735 ( .A1(n247), .A2(n279), .B1(\mem[25][23] ), .B2(n247), .ZN(
        n1337) );
  NR2XD0 U736 ( .A1(n278), .A2(n254), .ZN(n248) );
  MAOI22D0 U737 ( .A1(n248), .A2(n281), .B1(\mem[24][0] ), .B2(n248), .ZN(
        n1338) );
  MAOI22D0 U738 ( .A1(n248), .A2(n505), .B1(\mem[24][1] ), .B2(n248), .ZN(
        n1339) );
  MAOI22D0 U739 ( .A1(n248), .A2(n755), .B1(\mem[24][2] ), .B2(n248), .ZN(
        n1340) );
  MAOI22D0 U740 ( .A1(n248), .A2(n483), .B1(\mem[24][3] ), .B2(n248), .ZN(
        n1341) );
  MAOI22D0 U741 ( .A1(n248), .A2(n527), .B1(\mem[24][4] ), .B2(n248), .ZN(
        n1342) );
  MAOI22D0 U742 ( .A1(n248), .A2(n461), .B1(\mem[24][5] ), .B2(n248), .ZN(
        n1343) );
  MAOI22D0 U743 ( .A1(n248), .A2(n549), .B1(\mem[24][6] ), .B2(n248), .ZN(
        n1344) );
  MAOI22D0 U744 ( .A1(n248), .A2(n439), .B1(\mem[24][7] ), .B2(n248), .ZN(
        n1345) );
  MAOI22D0 U745 ( .A1(n248), .A2(n571), .B1(\mem[24][8] ), .B2(n248), .ZN(
        n1346) );
  MAOI22D0 U746 ( .A1(n248), .A2(n417), .B1(\mem[24][9] ), .B2(n248), .ZN(
        n1347) );
  MAOI22D0 U747 ( .A1(n248), .A2(n593), .B1(\mem[24][10] ), .B2(n248), .ZN(
        n1348) );
  MAOI22D0 U748 ( .A1(n248), .A2(n615), .B1(\mem[24][12] ), .B2(n248), .ZN(
        n1350) );
  MAOI22D0 U749 ( .A1(n248), .A2(n373), .B1(\mem[24][13] ), .B2(n248), .ZN(
        n1351) );
  MAOI22D0 U750 ( .A1(n248), .A2(n637), .B1(\mem[24][14] ), .B2(n248), .ZN(
        n1352) );
  MAOI22D0 U751 ( .A1(n248), .A2(n351), .B1(\mem[24][15] ), .B2(n248), .ZN(
        n1353) );
  MAOI22D0 U752 ( .A1(n248), .A2(n659), .B1(\mem[24][16] ), .B2(n248), .ZN(
        n1354) );
  MAOI22D0 U753 ( .A1(n248), .A2(n329), .B1(\mem[24][17] ), .B2(n248), .ZN(
        n1355) );
  MAOI22D0 U754 ( .A1(n248), .A2(n681), .B1(\mem[24][18] ), .B2(n248), .ZN(
        n1356) );
  MAOI22D0 U755 ( .A1(n248), .A2(n307), .B1(\mem[24][19] ), .B2(n248), .ZN(
        n1357) );
  MAOI22D0 U756 ( .A1(n248), .A2(n703), .B1(\mem[24][20] ), .B2(n248), .ZN(
        n1358) );
  MAOI22D0 U757 ( .A1(n248), .A2(n285), .B1(\mem[24][21] ), .B2(n248), .ZN(
        n1359) );
  MAOI22D0 U758 ( .A1(n248), .A2(n725), .B1(\mem[24][22] ), .B2(n248), .ZN(
        n1360) );
  MAOI22D0 U759 ( .A1(n248), .A2(n279), .B1(\mem[24][23] ), .B2(n248), .ZN(
        n1361) );
  CKND2D0 U760 ( .A1(write), .A2(n249), .ZN(n277) );
  NR2XD0 U761 ( .A1(n257), .A2(n277), .ZN(n250) );
  MAOI22D0 U762 ( .A1(n250), .A2(n281), .B1(\mem[23][0] ), .B2(n250), .ZN(
        n1362) );
  MAOI22D0 U763 ( .A1(n250), .A2(n505), .B1(\mem[23][1] ), .B2(n250), .ZN(
        n1363) );
  MAOI22D0 U764 ( .A1(n250), .A2(n483), .B1(\mem[23][3] ), .B2(n250), .ZN(
        n1365) );
  MAOI22D0 U765 ( .A1(n250), .A2(n527), .B1(\mem[23][4] ), .B2(n250), .ZN(
        n1366) );
  MAOI22D0 U766 ( .A1(n250), .A2(n461), .B1(\mem[23][5] ), .B2(n250), .ZN(
        n1367) );
  MAOI22D0 U767 ( .A1(n250), .A2(n549), .B1(\mem[23][6] ), .B2(n250), .ZN(
        n1368) );
  MAOI22D0 U768 ( .A1(n250), .A2(n439), .B1(\mem[23][7] ), .B2(n250), .ZN(
        n1369) );
  MAOI22D0 U769 ( .A1(n250), .A2(n571), .B1(\mem[23][8] ), .B2(n250), .ZN(
        n1370) );
  MAOI22D0 U770 ( .A1(n250), .A2(n417), .B1(\mem[23][9] ), .B2(n250), .ZN(
        n1371) );
  MAOI22D0 U771 ( .A1(n250), .A2(n593), .B1(\mem[23][10] ), .B2(n250), .ZN(
        n1372) );
  MAOI22D0 U772 ( .A1(n250), .A2(n395), .B1(\mem[23][11] ), .B2(n250), .ZN(
        n1373) );
  MAOI22D0 U773 ( .A1(n250), .A2(n615), .B1(\mem[23][12] ), .B2(n250), .ZN(
        n1374) );
  MAOI22D0 U774 ( .A1(n250), .A2(n373), .B1(\mem[23][13] ), .B2(n250), .ZN(
        n1375) );
  MAOI22D0 U775 ( .A1(n250), .A2(n637), .B1(\mem[23][14] ), .B2(n250), .ZN(
        n1376) );
  MAOI22D0 U776 ( .A1(n250), .A2(n351), .B1(\mem[23][15] ), .B2(n250), .ZN(
        n1377) );
  MAOI22D0 U777 ( .A1(n250), .A2(n659), .B1(\mem[23][16] ), .B2(n250), .ZN(
        n1378) );
  MAOI22D0 U778 ( .A1(n250), .A2(n681), .B1(\mem[23][18] ), .B2(n250), .ZN(
        n1380) );
  MAOI22D0 U779 ( .A1(n250), .A2(n307), .B1(\mem[23][19] ), .B2(n250), .ZN(
        n1381) );
  MAOI22D0 U780 ( .A1(n250), .A2(n703), .B1(\mem[23][20] ), .B2(n250), .ZN(
        n1382) );
  MAOI22D0 U781 ( .A1(n250), .A2(n285), .B1(\mem[23][21] ), .B2(n250), .ZN(
        n1383) );
  MAOI22D0 U782 ( .A1(n250), .A2(n725), .B1(\mem[23][22] ), .B2(n250), .ZN(
        n1384) );
  MAOI22D0 U783 ( .A1(n250), .A2(n279), .B1(\mem[23][23] ), .B2(n250), .ZN(
        n1385) );
  NR2XD0 U784 ( .A1(n258), .A2(n277), .ZN(n251) );
  MAOI22D0 U785 ( .A1(n251), .A2(n281), .B1(\mem[22][0] ), .B2(n251), .ZN(
        n1386) );
  MAOI22D0 U786 ( .A1(n251), .A2(n505), .B1(\mem[22][1] ), .B2(n251), .ZN(
        n1387) );
  MAOI22D0 U787 ( .A1(n251), .A2(n755), .B1(\mem[22][2] ), .B2(n251), .ZN(
        n1388) );
  MAOI22D0 U788 ( .A1(n251), .A2(n483), .B1(\mem[22][3] ), .B2(n251), .ZN(
        n1389) );
  MAOI22D0 U789 ( .A1(n251), .A2(n527), .B1(\mem[22][4] ), .B2(n251), .ZN(
        n1390) );
  MAOI22D0 U790 ( .A1(n251), .A2(n461), .B1(\mem[22][5] ), .B2(n251), .ZN(
        n1391) );
  MAOI22D0 U791 ( .A1(n251), .A2(n549), .B1(\mem[22][6] ), .B2(n251), .ZN(
        n1392) );
  MAOI22D0 U792 ( .A1(n251), .A2(n439), .B1(\mem[22][7] ), .B2(n251), .ZN(
        n1393) );
  MAOI22D0 U793 ( .A1(n251), .A2(n417), .B1(\mem[22][9] ), .B2(n251), .ZN(
        n1395) );
  MAOI22D0 U794 ( .A1(n251), .A2(n593), .B1(\mem[22][10] ), .B2(n251), .ZN(
        n1396) );
  MAOI22D0 U795 ( .A1(n251), .A2(n395), .B1(\mem[22][11] ), .B2(n251), .ZN(
        n1397) );
  MAOI22D0 U796 ( .A1(n251), .A2(n615), .B1(\mem[22][12] ), .B2(n251), .ZN(
        n1398) );
  MAOI22D0 U797 ( .A1(n251), .A2(n373), .B1(\mem[22][13] ), .B2(n251), .ZN(
        n1399) );
  MAOI22D0 U798 ( .A1(n251), .A2(n637), .B1(\mem[22][14] ), .B2(n251), .ZN(
        n1400) );
  MAOI22D0 U799 ( .A1(n251), .A2(n351), .B1(\mem[22][15] ), .B2(n251), .ZN(
        n1401) );
  MAOI22D0 U800 ( .A1(n251), .A2(n659), .B1(\mem[22][16] ), .B2(n251), .ZN(
        n1402) );
  MAOI22D0 U801 ( .A1(n251), .A2(n329), .B1(\mem[22][17] ), .B2(n251), .ZN(
        n1403) );
  MAOI22D0 U802 ( .A1(n251), .A2(n681), .B1(\mem[22][18] ), .B2(n251), .ZN(
        n1404) );
  MAOI22D0 U803 ( .A1(n251), .A2(n307), .B1(\mem[22][19] ), .B2(n251), .ZN(
        n1405) );
  MAOI22D0 U804 ( .A1(n251), .A2(n703), .B1(\mem[22][20] ), .B2(n251), .ZN(
        n1406) );
  MAOI22D0 U805 ( .A1(n251), .A2(n285), .B1(\mem[22][21] ), .B2(n251), .ZN(
        n1407) );
  MAOI22D0 U806 ( .A1(n251), .A2(n725), .B1(\mem[22][22] ), .B2(n251), .ZN(
        n1408) );
  NR2XD0 U807 ( .A1(n260), .A2(n277), .ZN(n273) );
  MAOI22D0 U808 ( .A1(n273), .A2(n281), .B1(\mem[21][0] ), .B2(n273), .ZN(
        n1410) );
  MAOI22D0 U809 ( .A1(n273), .A2(n505), .B1(\mem[21][1] ), .B2(n273), .ZN(
        n1411) );
  MAOI22D0 U810 ( .A1(n273), .A2(n755), .B1(\mem[21][2] ), .B2(n273), .ZN(
        n1412) );
  MAOI22D0 U811 ( .A1(n273), .A2(n483), .B1(\mem[21][3] ), .B2(n273), .ZN(
        n1413) );
  MAOI22D0 U812 ( .A1(n273), .A2(n527), .B1(\mem[21][4] ), .B2(n273), .ZN(
        n1414) );
  MAOI22D0 U813 ( .A1(n256), .A2(n351), .B1(\mem[28][15] ), .B2(n256), .ZN(
        n1257) );
  NR2XD0 U814 ( .A1(n257), .A2(n254), .ZN(n252) );
  MAOI22D0 U815 ( .A1(n252), .A2(n505), .B1(\mem[31][1] ), .B2(n252), .ZN(
        n1171) );
  MAOI22D0 U816 ( .A1(n252), .A2(n755), .B1(\mem[31][2] ), .B2(n252), .ZN(
        n1172) );
  MAOI22D0 U817 ( .A1(n252), .A2(n483), .B1(\mem[31][3] ), .B2(n252), .ZN(
        n1173) );
  MAOI22D0 U818 ( .A1(n252), .A2(n527), .B1(\mem[31][4] ), .B2(n252), .ZN(
        n1174) );
  MAOI22D0 U819 ( .A1(n252), .A2(n461), .B1(\mem[31][5] ), .B2(n252), .ZN(
        n1175) );
  MAOI22D0 U820 ( .A1(n252), .A2(n549), .B1(\mem[31][6] ), .B2(n252), .ZN(
        n1176) );
  MAOI22D0 U821 ( .A1(n252), .A2(n439), .B1(\mem[31][7] ), .B2(n252), .ZN(
        n1177) );
  MAOI22D0 U822 ( .A1(n252), .A2(n571), .B1(\mem[31][8] ), .B2(n252), .ZN(
        n1178) );
  MAOI22D0 U823 ( .A1(n252), .A2(n417), .B1(\mem[31][9] ), .B2(n252), .ZN(
        n1179) );
  MAOI22D0 U824 ( .A1(n252), .A2(n593), .B1(\mem[31][10] ), .B2(n252), .ZN(
        n1180) );
  MAOI22D0 U825 ( .A1(n252), .A2(n395), .B1(\mem[31][11] ), .B2(n252), .ZN(
        n1181) );
  MAOI22D0 U826 ( .A1(n252), .A2(n615), .B1(\mem[31][12] ), .B2(n252), .ZN(
        n1182) );
  MAOI22D0 U827 ( .A1(n252), .A2(n373), .B1(\mem[31][13] ), .B2(n252), .ZN(
        n1183) );
  MAOI22D0 U828 ( .A1(n252), .A2(n351), .B1(\mem[31][15] ), .B2(n252), .ZN(
        n1185) );
  MAOI22D0 U829 ( .A1(n252), .A2(n659), .B1(\mem[31][16] ), .B2(n252), .ZN(
        n1186) );
  MAOI22D0 U830 ( .A1(n252), .A2(n329), .B1(\mem[31][17] ), .B2(n252), .ZN(
        n1187) );
  MAOI22D0 U831 ( .A1(n252), .A2(n681), .B1(\mem[31][18] ), .B2(n252), .ZN(
        n1188) );
  MAOI22D0 U832 ( .A1(n252), .A2(n307), .B1(\mem[31][19] ), .B2(n252), .ZN(
        n1189) );
  MAOI22D0 U833 ( .A1(n252), .A2(n703), .B1(\mem[31][20] ), .B2(n252), .ZN(
        n1190) );
  MAOI22D0 U834 ( .A1(n252), .A2(n285), .B1(\mem[31][21] ), .B2(n252), .ZN(
        n1191) );
  MAOI22D0 U835 ( .A1(n252), .A2(n725), .B1(\mem[31][22] ), .B2(n252), .ZN(
        n1192) );
  MAOI22D0 U836 ( .A1(n252), .A2(n279), .B1(\mem[31][23] ), .B2(n252), .ZN(
        n1193) );
  NR2XD0 U837 ( .A1(n258), .A2(n254), .ZN(n253) );
  MAOI22D0 U838 ( .A1(n253), .A2(n281), .B1(\mem[30][0] ), .B2(n253), .ZN(
        n1194) );
  MAOI22D0 U839 ( .A1(n253), .A2(n505), .B1(\mem[30][1] ), .B2(n253), .ZN(
        n1195) );
  MAOI22D0 U840 ( .A1(n253), .A2(n755), .B1(\mem[30][2] ), .B2(n253), .ZN(
        n1196) );
  MAOI22D0 U841 ( .A1(n253), .A2(n483), .B1(\mem[30][3] ), .B2(n253), .ZN(
        n1197) );
  MAOI22D0 U842 ( .A1(n253), .A2(n527), .B1(\mem[30][4] ), .B2(n253), .ZN(
        n1198) );
  MAOI22D0 U843 ( .A1(n253), .A2(n549), .B1(\mem[30][6] ), .B2(n253), .ZN(
        n1200) );
  MAOI22D0 U844 ( .A1(n253), .A2(n439), .B1(\mem[30][7] ), .B2(n253), .ZN(
        n1201) );
  MAOI22D0 U845 ( .A1(n253), .A2(n571), .B1(\mem[30][8] ), .B2(n253), .ZN(
        n1202) );
  MAOI22D0 U846 ( .A1(n253), .A2(n417), .B1(\mem[30][9] ), .B2(n253), .ZN(
        n1203) );
  MAOI22D0 U847 ( .A1(n253), .A2(n593), .B1(\mem[30][10] ), .B2(n253), .ZN(
        n1204) );
  MAOI22D0 U848 ( .A1(n253), .A2(n395), .B1(\mem[30][11] ), .B2(n253), .ZN(
        n1205) );
  MAOI22D0 U849 ( .A1(n253), .A2(n615), .B1(\mem[30][12] ), .B2(n253), .ZN(
        n1206) );
  MAOI22D0 U850 ( .A1(n253), .A2(n373), .B1(\mem[30][13] ), .B2(n253), .ZN(
        n1207) );
  MAOI22D0 U851 ( .A1(n253), .A2(n637), .B1(\mem[30][14] ), .B2(n253), .ZN(
        n1208) );
  MAOI22D0 U852 ( .A1(n253), .A2(n351), .B1(\mem[30][15] ), .B2(n253), .ZN(
        n1209) );
  MAOI22D0 U853 ( .A1(n253), .A2(n659), .B1(\mem[30][16] ), .B2(n253), .ZN(
        n1210) );
  MAOI22D0 U854 ( .A1(n253), .A2(n329), .B1(\mem[30][17] ), .B2(n253), .ZN(
        n1211) );
  MAOI22D0 U855 ( .A1(n253), .A2(n681), .B1(\mem[30][18] ), .B2(n253), .ZN(
        n1212) );
  MAOI22D0 U856 ( .A1(n253), .A2(n307), .B1(\mem[30][19] ), .B2(n253), .ZN(
        n1213) );
  MAOI22D0 U857 ( .A1(n253), .A2(n285), .B1(\mem[30][21] ), .B2(n253), .ZN(
        n1215) );
  MAOI22D0 U858 ( .A1(n253), .A2(n725), .B1(\mem[30][22] ), .B2(n253), .ZN(
        n1216) );
  MAOI22D0 U859 ( .A1(n253), .A2(n279), .B1(\mem[30][23] ), .B2(n253), .ZN(
        n1217) );
  NR2XD0 U860 ( .A1(n260), .A2(n254), .ZN(n255) );
  MAOI22D0 U861 ( .A1(n255), .A2(n281), .B1(\mem[29][0] ), .B2(n255), .ZN(
        n1218) );
  MAOI22D0 U862 ( .A1(n255), .A2(n505), .B1(\mem[29][1] ), .B2(n255), .ZN(
        n1219) );
  MAOI22D0 U863 ( .A1(n255), .A2(n755), .B1(\mem[29][2] ), .B2(n255), .ZN(
        n1220) );
  MAOI22D0 U864 ( .A1(n255), .A2(n483), .B1(\mem[29][3] ), .B2(n255), .ZN(
        n1221) );
  MAOI22D0 U865 ( .A1(n255), .A2(n527), .B1(\mem[29][4] ), .B2(n255), .ZN(
        n1222) );
  MAOI22D0 U866 ( .A1(n255), .A2(n461), .B1(\mem[29][5] ), .B2(n255), .ZN(
        n1223) );
  MAOI22D0 U867 ( .A1(n255), .A2(n549), .B1(\mem[29][6] ), .B2(n255), .ZN(
        n1224) );
  MAOI22D0 U868 ( .A1(n255), .A2(n439), .B1(\mem[29][7] ), .B2(n255), .ZN(
        n1225) );
  MAOI22D0 U869 ( .A1(n255), .A2(n571), .B1(\mem[29][8] ), .B2(n255), .ZN(
        n1226) );
  MAOI22D0 U870 ( .A1(n255), .A2(n417), .B1(\mem[29][9] ), .B2(n255), .ZN(
        n1227) );
  MAOI22D0 U871 ( .A1(n255), .A2(n593), .B1(\mem[29][10] ), .B2(n255), .ZN(
        n1228) );
  MAOI22D0 U872 ( .A1(n255), .A2(n615), .B1(\mem[29][12] ), .B2(n255), .ZN(
        n1230) );
  MAOI22D0 U873 ( .A1(n255), .A2(n373), .B1(\mem[29][13] ), .B2(n255), .ZN(
        n1231) );
  MAOI22D0 U874 ( .A1(n255), .A2(n637), .B1(\mem[29][14] ), .B2(n255), .ZN(
        n1232) );
  MAOI22D0 U875 ( .A1(n255), .A2(n351), .B1(\mem[29][15] ), .B2(n255), .ZN(
        n1233) );
  MAOI22D0 U876 ( .A1(n255), .A2(n659), .B1(\mem[29][16] ), .B2(n255), .ZN(
        n1234) );
  MAOI22D0 U877 ( .A1(n255), .A2(n329), .B1(\mem[29][17] ), .B2(n255), .ZN(
        n1235) );
  MAOI22D0 U878 ( .A1(n255), .A2(n681), .B1(\mem[29][18] ), .B2(n255), .ZN(
        n1236) );
  MAOI22D0 U879 ( .A1(n255), .A2(n307), .B1(\mem[29][19] ), .B2(n255), .ZN(
        n1237) );
  MAOI22D0 U880 ( .A1(n255), .A2(n703), .B1(\mem[29][20] ), .B2(n255), .ZN(
        n1238) );
  MAOI22D0 U881 ( .A1(n255), .A2(n285), .B1(\mem[29][21] ), .B2(n255), .ZN(
        n1239) );
  MAOI22D0 U882 ( .A1(n255), .A2(n725), .B1(\mem[29][22] ), .B2(n255), .ZN(
        n1240) );
  MAOI22D0 U883 ( .A1(n255), .A2(n279), .B1(\mem[29][23] ), .B2(n255), .ZN(
        n1241) );
  MAOI22D0 U884 ( .A1(n256), .A2(n281), .B1(\mem[28][0] ), .B2(n256), .ZN(
        n1242) );
  MAOI22D0 U885 ( .A1(n256), .A2(n505), .B1(\mem[28][1] ), .B2(n256), .ZN(
        n1243) );
  MAOI22D0 U886 ( .A1(n256), .A2(n483), .B1(\mem[28][3] ), .B2(n256), .ZN(
        n1245) );
  MAOI22D0 U887 ( .A1(n256), .A2(n527), .B1(\mem[28][4] ), .B2(n256), .ZN(
        n1246) );
  MAOI22D0 U888 ( .A1(n256), .A2(n461), .B1(\mem[28][5] ), .B2(n256), .ZN(
        n1247) );
  MAOI22D0 U889 ( .A1(n256), .A2(n549), .B1(\mem[28][6] ), .B2(n256), .ZN(
        n1248) );
  MAOI22D0 U890 ( .A1(n256), .A2(n439), .B1(\mem[28][7] ), .B2(n256), .ZN(
        n1249) );
  MAOI22D0 U891 ( .A1(n256), .A2(n571), .B1(\mem[28][8] ), .B2(n256), .ZN(
        n1250) );
  MAOI22D0 U892 ( .A1(n256), .A2(n417), .B1(\mem[28][9] ), .B2(n256), .ZN(
        n1251) );
  MAOI22D0 U893 ( .A1(n256), .A2(n593), .B1(\mem[28][10] ), .B2(n256), .ZN(
        n1252) );
  MAOI22D0 U894 ( .A1(n256), .A2(n395), .B1(\mem[28][11] ), .B2(n256), .ZN(
        n1253) );
  MAOI22D0 U895 ( .A1(n256), .A2(n615), .B1(\mem[28][12] ), .B2(n256), .ZN(
        n1254) );
  MAOI22D0 U896 ( .A1(n256), .A2(n373), .B1(\mem[28][13] ), .B2(n256), .ZN(
        n1255) );
  MAOI22D0 U897 ( .A1(n256), .A2(n637), .B1(\mem[28][14] ), .B2(n256), .ZN(
        n1256) );
  MAOI22D0 U898 ( .A1(n273), .A2(n461), .B1(\mem[21][5] ), .B2(n273), .ZN(
        n1415) );
  NR2XD0 U899 ( .A1(n257), .A2(n265), .ZN(n282) );
  MAOI22D0 U900 ( .A1(n282), .A2(n285), .B1(\mem[15][21] ), .B2(n282), .ZN(
        n1575) );
  MAOI22D0 U901 ( .A1(n282), .A2(n725), .B1(\mem[15][22] ), .B2(n282), .ZN(
        n1576) );
  MAOI22D0 U902 ( .A1(n282), .A2(n279), .B1(\mem[15][23] ), .B2(n282), .ZN(
        n1577) );
  NR2XD0 U903 ( .A1(n258), .A2(n265), .ZN(n259) );
  MAOI22D0 U904 ( .A1(n259), .A2(n281), .B1(\mem[14][0] ), .B2(n259), .ZN(
        n1578) );
  MAOI22D0 U905 ( .A1(n259), .A2(n505), .B1(\mem[14][1] ), .B2(n259), .ZN(
        n1579) );
  MAOI22D0 U906 ( .A1(n259), .A2(n755), .B1(\mem[14][2] ), .B2(n259), .ZN(
        n1580) );
  MAOI22D0 U907 ( .A1(n259), .A2(n483), .B1(\mem[14][3] ), .B2(n259), .ZN(
        n1581) );
  MAOI22D0 U908 ( .A1(n259), .A2(n527), .B1(\mem[14][4] ), .B2(n259), .ZN(
        n1582) );
  MAOI22D0 U909 ( .A1(n259), .A2(n461), .B1(\mem[14][5] ), .B2(n259), .ZN(
        n1583) );
  MAOI22D0 U910 ( .A1(n259), .A2(n549), .B1(\mem[14][6] ), .B2(n259), .ZN(
        n1584) );
  MAOI22D0 U911 ( .A1(n259), .A2(n439), .B1(\mem[14][7] ), .B2(n259), .ZN(
        n1585) );
  MAOI22D0 U912 ( .A1(n259), .A2(n571), .B1(\mem[14][8] ), .B2(n259), .ZN(
        n1586) );
  MAOI22D0 U913 ( .A1(n259), .A2(n417), .B1(\mem[14][9] ), .B2(n259), .ZN(
        n1587) );
  MAOI22D0 U914 ( .A1(n259), .A2(n593), .B1(\mem[14][10] ), .B2(n259), .ZN(
        n1588) );
  MAOI22D0 U915 ( .A1(n259), .A2(n615), .B1(\mem[14][12] ), .B2(n259), .ZN(
        n1590) );
  MAOI22D0 U916 ( .A1(n259), .A2(n373), .B1(\mem[14][13] ), .B2(n259), .ZN(
        n1591) );
  MAOI22D0 U917 ( .A1(n259), .A2(n637), .B1(\mem[14][14] ), .B2(n259), .ZN(
        n1592) );
  MAOI22D0 U918 ( .A1(n259), .A2(n351), .B1(\mem[14][15] ), .B2(n259), .ZN(
        n1593) );
  MAOI22D0 U919 ( .A1(n259), .A2(n659), .B1(\mem[14][16] ), .B2(n259), .ZN(
        n1594) );
  MAOI22D0 U920 ( .A1(n259), .A2(n329), .B1(\mem[14][17] ), .B2(n259), .ZN(
        n1595) );
  MAOI22D0 U921 ( .A1(n259), .A2(n681), .B1(\mem[14][18] ), .B2(n259), .ZN(
        n1596) );
  MAOI22D0 U922 ( .A1(n259), .A2(n307), .B1(\mem[14][19] ), .B2(n259), .ZN(
        n1597) );
  MAOI22D0 U923 ( .A1(n259), .A2(n703), .B1(\mem[14][20] ), .B2(n259), .ZN(
        n1598) );
  MAOI22D0 U924 ( .A1(n259), .A2(n285), .B1(\mem[14][21] ), .B2(n259), .ZN(
        n1599) );
  MAOI22D0 U925 ( .A1(n259), .A2(n725), .B1(\mem[14][22] ), .B2(n259), .ZN(
        n1600) );
  MAOI22D0 U926 ( .A1(n259), .A2(n279), .B1(\mem[14][23] ), .B2(n259), .ZN(
        n1601) );
  NR2XD0 U927 ( .A1(n260), .A2(n265), .ZN(n261) );
  MAOI22D0 U928 ( .A1(n261), .A2(n281), .B1(\mem[13][0] ), .B2(n261), .ZN(
        n1602) );
  MAOI22D0 U929 ( .A1(n261), .A2(n505), .B1(\mem[13][1] ), .B2(n261), .ZN(
        n1603) );
  MAOI22D0 U930 ( .A1(n261), .A2(n483), .B1(\mem[13][3] ), .B2(n261), .ZN(
        n1605) );
  MAOI22D0 U931 ( .A1(n261), .A2(n527), .B1(\mem[13][4] ), .B2(n261), .ZN(
        n1606) );
  MAOI22D0 U932 ( .A1(n261), .A2(n461), .B1(\mem[13][5] ), .B2(n261), .ZN(
        n1607) );
  MAOI22D0 U933 ( .A1(n261), .A2(n549), .B1(\mem[13][6] ), .B2(n261), .ZN(
        n1608) );
  MAOI22D0 U934 ( .A1(n261), .A2(n439), .B1(\mem[13][7] ), .B2(n261), .ZN(
        n1609) );
  MAOI22D0 U935 ( .A1(n261), .A2(n571), .B1(\mem[13][8] ), .B2(n261), .ZN(
        n1610) );
  MAOI22D0 U936 ( .A1(n261), .A2(n417), .B1(\mem[13][9] ), .B2(n261), .ZN(
        n1611) );
  MAOI22D0 U937 ( .A1(n261), .A2(n593), .B1(\mem[13][10] ), .B2(n261), .ZN(
        n1612) );
  MAOI22D0 U938 ( .A1(n261), .A2(n395), .B1(\mem[13][11] ), .B2(n261), .ZN(
        n1613) );
  MAOI22D0 U939 ( .A1(n261), .A2(n615), .B1(\mem[13][12] ), .B2(n261), .ZN(
        n1614) );
  MAOI22D0 U940 ( .A1(n261), .A2(n373), .B1(\mem[13][13] ), .B2(n261), .ZN(
        n1615) );
  MAOI22D0 U941 ( .A1(n261), .A2(n637), .B1(\mem[13][14] ), .B2(n261), .ZN(
        n1616) );
  MAOI22D0 U942 ( .A1(n261), .A2(n351), .B1(\mem[13][15] ), .B2(n261), .ZN(
        n1617) );
  MAOI22D0 U943 ( .A1(n261), .A2(n659), .B1(\mem[13][16] ), .B2(n261), .ZN(
        n1618) );
  MAOI22D0 U944 ( .A1(n261), .A2(n681), .B1(\mem[13][18] ), .B2(n261), .ZN(
        n1620) );
  MAOI22D0 U945 ( .A1(n261), .A2(n307), .B1(\mem[13][19] ), .B2(n261), .ZN(
        n1621) );
  MAOI22D0 U946 ( .A1(n261), .A2(n703), .B1(\mem[13][20] ), .B2(n261), .ZN(
        n1622) );
  MAOI22D0 U947 ( .A1(n261), .A2(n285), .B1(\mem[13][21] ), .B2(n261), .ZN(
        n1623) );
  MAOI22D0 U948 ( .A1(n261), .A2(n725), .B1(\mem[13][22] ), .B2(n261), .ZN(
        n1624) );
  MAOI22D0 U949 ( .A1(n261), .A2(n279), .B1(\mem[13][23] ), .B2(n261), .ZN(
        n1625) );
  NR2XD0 U950 ( .A1(n268), .A2(n265), .ZN(n262) );
  MAOI22D0 U951 ( .A1(n262), .A2(n281), .B1(\mem[12][0] ), .B2(n262), .ZN(
        n1626) );
  MAOI22D0 U952 ( .A1(n262), .A2(n505), .B1(\mem[12][1] ), .B2(n262), .ZN(
        n1627) );
  MAOI22D0 U953 ( .A1(n262), .A2(n755), .B1(\mem[12][2] ), .B2(n262), .ZN(
        n1628) );
  MAOI22D0 U954 ( .A1(n262), .A2(n483), .B1(\mem[12][3] ), .B2(n262), .ZN(
        n1629) );
  MAOI22D0 U955 ( .A1(n262), .A2(n527), .B1(\mem[12][4] ), .B2(n262), .ZN(
        n1630) );
  MAOI22D0 U956 ( .A1(n262), .A2(n461), .B1(\mem[12][5] ), .B2(n262), .ZN(
        n1631) );
  MAOI22D0 U957 ( .A1(n262), .A2(n549), .B1(\mem[12][6] ), .B2(n262), .ZN(
        n1632) );
  MAOI22D0 U958 ( .A1(n262), .A2(n439), .B1(\mem[12][7] ), .B2(n262), .ZN(
        n1633) );
  MAOI22D0 U959 ( .A1(n262), .A2(n417), .B1(\mem[12][9] ), .B2(n262), .ZN(
        n1635) );
  MAOI22D0 U960 ( .A1(n262), .A2(n593), .B1(\mem[12][10] ), .B2(n262), .ZN(
        n1636) );
  MAOI22D0 U961 ( .A1(n262), .A2(n395), .B1(\mem[12][11] ), .B2(n262), .ZN(
        n1637) );
  MAOI22D0 U962 ( .A1(n262), .A2(n615), .B1(\mem[12][12] ), .B2(n262), .ZN(
        n1638) );
  MAOI22D0 U963 ( .A1(n262), .A2(n373), .B1(\mem[12][13] ), .B2(n262), .ZN(
        n1639) );
  MAOI22D0 U964 ( .A1(n262), .A2(n637), .B1(\mem[12][14] ), .B2(n262), .ZN(
        n1640) );
  MAOI22D0 U965 ( .A1(n262), .A2(n351), .B1(\mem[12][15] ), .B2(n262), .ZN(
        n1641) );
  MAOI22D0 U966 ( .A1(n262), .A2(n659), .B1(\mem[12][16] ), .B2(n262), .ZN(
        n1642) );
  MAOI22D0 U967 ( .A1(n262), .A2(n329), .B1(\mem[12][17] ), .B2(n262), .ZN(
        n1643) );
  MAOI22D0 U968 ( .A1(n262), .A2(n681), .B1(\mem[12][18] ), .B2(n262), .ZN(
        n1644) );
  MAOI22D0 U969 ( .A1(n262), .A2(n307), .B1(\mem[12][19] ), .B2(n262), .ZN(
        n1645) );
  MAOI22D0 U970 ( .A1(n262), .A2(n703), .B1(\mem[12][20] ), .B2(n262), .ZN(
        n1646) );
  MAOI22D0 U971 ( .A1(n262), .A2(n285), .B1(\mem[12][21] ), .B2(n262), .ZN(
        n1647) );
  MAOI22D0 U972 ( .A1(n262), .A2(n725), .B1(\mem[12][22] ), .B2(n262), .ZN(
        n1648) );
  NR2XD0 U973 ( .A1(n270), .A2(n265), .ZN(n263) );
  MAOI22D0 U974 ( .A1(n263), .A2(n281), .B1(\mem[11][0] ), .B2(n263), .ZN(
        n1650) );
  MAOI22D0 U975 ( .A1(n263), .A2(n505), .B1(\mem[11][1] ), .B2(n263), .ZN(
        n1651) );
  MAOI22D0 U976 ( .A1(n263), .A2(n755), .B1(\mem[11][2] ), .B2(n263), .ZN(
        n1652) );
  MAOI22D0 U977 ( .A1(n263), .A2(n483), .B1(\mem[11][3] ), .B2(n263), .ZN(
        n1653) );
  MAOI22D0 U978 ( .A1(n263), .A2(n527), .B1(\mem[11][4] ), .B2(n263), .ZN(
        n1654) );
  MAOI22D0 U979 ( .A1(n263), .A2(n461), .B1(\mem[11][5] ), .B2(n263), .ZN(
        n1655) );
  MAOI22D0 U980 ( .A1(n263), .A2(n549), .B1(\mem[11][6] ), .B2(n263), .ZN(
        n1656) );
  MAOI22D0 U981 ( .A1(n263), .A2(n439), .B1(\mem[11][7] ), .B2(n263), .ZN(
        n1657) );
  MAOI22D0 U982 ( .A1(n263), .A2(n571), .B1(\mem[11][8] ), .B2(n263), .ZN(
        n1658) );
  MAOI22D0 U983 ( .A1(n263), .A2(n417), .B1(\mem[11][9] ), .B2(n263), .ZN(
        n1659) );
  MAOI22D0 U984 ( .A1(n263), .A2(n593), .B1(\mem[11][10] ), .B2(n263), .ZN(
        n1660) );
  MAOI22D0 U985 ( .A1(n263), .A2(n395), .B1(\mem[11][11] ), .B2(n263), .ZN(
        n1661) );
  MAOI22D0 U986 ( .A1(n263), .A2(n615), .B1(\mem[11][12] ), .B2(n263), .ZN(
        n1662) );
  MAOI22D0 U987 ( .A1(n263), .A2(n373), .B1(\mem[11][13] ), .B2(n263), .ZN(
        n1663) );
  MAOI22D0 U988 ( .A1(n263), .A2(n351), .B1(\mem[11][15] ), .B2(n263), .ZN(
        n1665) );
  MAOI22D0 U989 ( .A1(n263), .A2(n659), .B1(\mem[11][16] ), .B2(n263), .ZN(
        n1666) );
  MAOI22D0 U990 ( .A1(n263), .A2(n329), .B1(\mem[11][17] ), .B2(n263), .ZN(
        n1667) );
  MAOI22D0 U991 ( .A1(n263), .A2(n681), .B1(\mem[11][18] ), .B2(n263), .ZN(
        n1668) );
  MAOI22D0 U992 ( .A1(n263), .A2(n307), .B1(\mem[11][19] ), .B2(n263), .ZN(
        n1669) );
  MAOI22D0 U993 ( .A1(n263), .A2(n703), .B1(\mem[11][20] ), .B2(n263), .ZN(
        n1670) );
  MAOI22D0 U994 ( .A1(n263), .A2(n285), .B1(\mem[11][21] ), .B2(n263), .ZN(
        n1671) );
  MAOI22D0 U995 ( .A1(n263), .A2(n725), .B1(\mem[11][22] ), .B2(n263), .ZN(
        n1672) );
  MAOI22D0 U996 ( .A1(n263), .A2(n279), .B1(\mem[11][23] ), .B2(n263), .ZN(
        n1673) );
  NR2XD0 U997 ( .A1(n272), .A2(n265), .ZN(n264) );
  MAOI22D0 U998 ( .A1(n264), .A2(n281), .B1(\mem[10][0] ), .B2(n264), .ZN(
        n1674) );
  MAOI22D0 U999 ( .A1(n264), .A2(n505), .B1(\mem[10][1] ), .B2(n264), .ZN(
        n1675) );
  MAOI22D0 U1000 ( .A1(n264), .A2(n755), .B1(\mem[10][2] ), .B2(n264), .ZN(
        n1676) );
  MAOI22D0 U1001 ( .A1(n264), .A2(n483), .B1(\mem[10][3] ), .B2(n264), .ZN(
        n1677) );
  MAOI22D0 U1002 ( .A1(n264), .A2(n527), .B1(\mem[10][4] ), .B2(n264), .ZN(
        n1678) );
  MAOI22D0 U1003 ( .A1(n264), .A2(n549), .B1(\mem[10][6] ), .B2(n264), .ZN(
        n1680) );
  MAOI22D0 U1004 ( .A1(n264), .A2(n439), .B1(\mem[10][7] ), .B2(n264), .ZN(
        n1681) );
  MAOI22D0 U1005 ( .A1(n264), .A2(n571), .B1(\mem[10][8] ), .B2(n264), .ZN(
        n1682) );
  MAOI22D0 U1006 ( .A1(n264), .A2(n417), .B1(\mem[10][9] ), .B2(n264), .ZN(
        n1683) );
  MAOI22D0 U1007 ( .A1(n264), .A2(n593), .B1(\mem[10][10] ), .B2(n264), .ZN(
        n1684) );
  MAOI22D0 U1008 ( .A1(n264), .A2(n395), .B1(\mem[10][11] ), .B2(n264), .ZN(
        n1685) );
  MAOI22D0 U1009 ( .A1(n264), .A2(n615), .B1(\mem[10][12] ), .B2(n264), .ZN(
        n1686) );
  MAOI22D0 U1010 ( .A1(n264), .A2(n373), .B1(\mem[10][13] ), .B2(n264), .ZN(
        n1687) );
  MAOI22D0 U1011 ( .A1(n264), .A2(n637), .B1(\mem[10][14] ), .B2(n264), .ZN(
        n1688) );
  MAOI22D0 U1012 ( .A1(n264), .A2(n351), .B1(\mem[10][15] ), .B2(n264), .ZN(
        n1689) );
  MAOI22D0 U1013 ( .A1(n264), .A2(n659), .B1(\mem[10][16] ), .B2(n264), .ZN(
        n1690) );
  MAOI22D0 U1014 ( .A1(n264), .A2(n329), .B1(\mem[10][17] ), .B2(n264), .ZN(
        n1691) );
  MAOI22D0 U1015 ( .A1(n264), .A2(n681), .B1(\mem[10][18] ), .B2(n264), .ZN(
        n1692) );
  MAOI22D0 U1016 ( .A1(n264), .A2(n307), .B1(\mem[10][19] ), .B2(n264), .ZN(
        n1693) );
  MAOI22D0 U1017 ( .A1(n264), .A2(n285), .B1(\mem[10][21] ), .B2(n264), .ZN(
        n1695) );
  MAOI22D0 U1018 ( .A1(n264), .A2(n725), .B1(\mem[10][22] ), .B2(n264), .ZN(
        n1696) );
  MAOI22D0 U1019 ( .A1(n264), .A2(n279), .B1(\mem[10][23] ), .B2(n264), .ZN(
        n1697) );
  NR2XD0 U1020 ( .A1(n275), .A2(n265), .ZN(n266) );
  MAOI22D0 U1021 ( .A1(n266), .A2(n281), .B1(\mem[9][0] ), .B2(n266), .ZN(
        n1698) );
  MAOI22D0 U1022 ( .A1(n266), .A2(n505), .B1(\mem[9][1] ), .B2(n266), .ZN(
        n1699) );
  MAOI22D0 U1023 ( .A1(n266), .A2(n755), .B1(\mem[9][2] ), .B2(n266), .ZN(
        n1700) );
  MAOI22D0 U1024 ( .A1(n266), .A2(n483), .B1(\mem[9][3] ), .B2(n266), .ZN(
        n1701) );
  MAOI22D0 U1025 ( .A1(n266), .A2(n527), .B1(\mem[9][4] ), .B2(n266), .ZN(
        n1702) );
  MAOI22D0 U1026 ( .A1(n266), .A2(n461), .B1(\mem[9][5] ), .B2(n266), .ZN(
        n1703) );
  MAOI22D0 U1027 ( .A1(n266), .A2(n549), .B1(\mem[9][6] ), .B2(n266), .ZN(
        n1704) );
  MAOI22D0 U1028 ( .A1(n266), .A2(n439), .B1(\mem[9][7] ), .B2(n266), .ZN(
        n1705) );
  MAOI22D0 U1029 ( .A1(n266), .A2(n571), .B1(\mem[9][8] ), .B2(n266), .ZN(
        n1706) );
  MAOI22D0 U1030 ( .A1(n266), .A2(n417), .B1(\mem[9][9] ), .B2(n266), .ZN(
        n1707) );
  MAOI22D0 U1031 ( .A1(n266), .A2(n593), .B1(\mem[9][10] ), .B2(n266), .ZN(
        n1708) );
  MAOI22D0 U1032 ( .A1(n266), .A2(n615), .B1(\mem[9][12] ), .B2(n266), .ZN(
        n1710) );
  MAOI22D0 U1033 ( .A1(n266), .A2(n373), .B1(\mem[9][13] ), .B2(n266), .ZN(
        n1711) );
  MAOI22D0 U1034 ( .A1(n266), .A2(n637), .B1(\mem[9][14] ), .B2(n266), .ZN(
        n1712) );
  MAOI22D0 U1035 ( .A1(n266), .A2(n351), .B1(\mem[9][15] ), .B2(n266), .ZN(
        n1713) );
  MAOI22D0 U1036 ( .A1(n266), .A2(n659), .B1(\mem[9][16] ), .B2(n266), .ZN(
        n1714) );
  MAOI22D0 U1037 ( .A1(n266), .A2(n329), .B1(\mem[9][17] ), .B2(n266), .ZN(
        n1715) );
  MAOI22D0 U1038 ( .A1(n266), .A2(n681), .B1(\mem[9][18] ), .B2(n266), .ZN(
        n1716) );
  MAOI22D0 U1039 ( .A1(n266), .A2(n307), .B1(\mem[9][19] ), .B2(n266), .ZN(
        n1717) );
  MAOI22D0 U1040 ( .A1(n266), .A2(n703), .B1(\mem[9][20] ), .B2(n266), .ZN(
        n1718) );
  MAOI22D0 U1041 ( .A1(n266), .A2(n285), .B1(\mem[9][21] ), .B2(n266), .ZN(
        n1719) );
  MAOI22D0 U1042 ( .A1(n266), .A2(n725), .B1(\mem[9][22] ), .B2(n266), .ZN(
        n1720) );
  MAOI22D0 U1043 ( .A1(n266), .A2(n279), .B1(\mem[9][23] ), .B2(n266), .ZN(
        n1721) );
  MAOI22D0 U1044 ( .A1(n267), .A2(n281), .B1(\mem[8][0] ), .B2(n267), .ZN(
        n1722) );
  MAOI22D0 U1045 ( .A1(n267), .A2(n505), .B1(\mem[8][1] ), .B2(n267), .ZN(
        n1723) );
  MAOI22D0 U1046 ( .A1(n267), .A2(n483), .B1(\mem[8][3] ), .B2(n267), .ZN(
        n1725) );
  MAOI22D0 U1047 ( .A1(n267), .A2(n527), .B1(\mem[8][4] ), .B2(n267), .ZN(
        n1726) );
  MAOI22D0 U1048 ( .A1(n267), .A2(n461), .B1(\mem[8][5] ), .B2(n267), .ZN(
        n1727) );
  MAOI22D0 U1049 ( .A1(n267), .A2(n549), .B1(\mem[8][6] ), .B2(n267), .ZN(
        n1728) );
  MAOI22D0 U1050 ( .A1(n267), .A2(n439), .B1(\mem[8][7] ), .B2(n267), .ZN(
        n1729) );
  MAOI22D0 U1051 ( .A1(n267), .A2(n571), .B1(\mem[8][8] ), .B2(n267), .ZN(
        n1730) );
  MAOI22D0 U1052 ( .A1(n282), .A2(n307), .B1(\mem[15][19] ), .B2(n282), .ZN(
        n1573) );
  MAOI22D0 U1053 ( .A1(n273), .A2(n439), .B1(\mem[21][7] ), .B2(n273), .ZN(
        n1417) );
  MAOI22D0 U1054 ( .A1(n273), .A2(n571), .B1(\mem[21][8] ), .B2(n273), .ZN(
        n1418) );
  MAOI22D0 U1055 ( .A1(n273), .A2(n417), .B1(\mem[21][9] ), .B2(n273), .ZN(
        n1419) );
  MAOI22D0 U1056 ( .A1(n273), .A2(n593), .B1(\mem[21][10] ), .B2(n273), .ZN(
        n1420) );
  MAOI22D0 U1057 ( .A1(n273), .A2(n395), .B1(\mem[21][11] ), .B2(n273), .ZN(
        n1421) );
  MAOI22D0 U1058 ( .A1(n273), .A2(n615), .B1(\mem[21][12] ), .B2(n273), .ZN(
        n1422) );
  MAOI22D0 U1059 ( .A1(n273), .A2(n373), .B1(\mem[21][13] ), .B2(n273), .ZN(
        n1423) );
  MAOI22D0 U1060 ( .A1(n273), .A2(n351), .B1(\mem[21][15] ), .B2(n273), .ZN(
        n1425) );
  MAOI22D0 U1061 ( .A1(n273), .A2(n659), .B1(\mem[21][16] ), .B2(n273), .ZN(
        n1426) );
  MAOI22D0 U1062 ( .A1(n273), .A2(n329), .B1(\mem[21][17] ), .B2(n273), .ZN(
        n1427) );
  MAOI22D0 U1063 ( .A1(n273), .A2(n681), .B1(\mem[21][18] ), .B2(n273), .ZN(
        n1428) );
  MAOI22D0 U1064 ( .A1(n273), .A2(n307), .B1(\mem[21][19] ), .B2(n273), .ZN(
        n1429) );
  MAOI22D0 U1065 ( .A1(n273), .A2(n703), .B1(\mem[21][20] ), .B2(n273), .ZN(
        n1430) );
  MAOI22D0 U1066 ( .A1(n273), .A2(n285), .B1(\mem[21][21] ), .B2(n273), .ZN(
        n1431) );
  MAOI22D0 U1067 ( .A1(n273), .A2(n725), .B1(\mem[21][22] ), .B2(n273), .ZN(
        n1432) );
  MAOI22D0 U1068 ( .A1(n273), .A2(n279), .B1(\mem[21][23] ), .B2(n273), .ZN(
        n1433) );
  NR2XD0 U1069 ( .A1(n268), .A2(n277), .ZN(n269) );
  MAOI22D0 U1070 ( .A1(n269), .A2(n281), .B1(\mem[20][0] ), .B2(n269), .ZN(
        n1434) );
  MAOI22D0 U1071 ( .A1(n269), .A2(n505), .B1(\mem[20][1] ), .B2(n269), .ZN(
        n1435) );
  MAOI22D0 U1072 ( .A1(n269), .A2(n755), .B1(\mem[20][2] ), .B2(n269), .ZN(
        n1436) );
  MAOI22D0 U1073 ( .A1(n269), .A2(n483), .B1(\mem[20][3] ), .B2(n269), .ZN(
        n1437) );
  MAOI22D0 U1074 ( .A1(n269), .A2(n527), .B1(\mem[20][4] ), .B2(n269), .ZN(
        n1438) );
  MAOI22D0 U1075 ( .A1(n269), .A2(n549), .B1(\mem[20][6] ), .B2(n269), .ZN(
        n1440) );
  MAOI22D0 U1076 ( .A1(n269), .A2(n439), .B1(\mem[20][7] ), .B2(n269), .ZN(
        n1441) );
  MAOI22D0 U1077 ( .A1(n269), .A2(n571), .B1(\mem[20][8] ), .B2(n269), .ZN(
        n1442) );
  MAOI22D0 U1078 ( .A1(n269), .A2(n417), .B1(\mem[20][9] ), .B2(n269), .ZN(
        n1443) );
  MAOI22D0 U1079 ( .A1(n269), .A2(n593), .B1(\mem[20][10] ), .B2(n269), .ZN(
        n1444) );
  MAOI22D0 U1080 ( .A1(n269), .A2(n395), .B1(\mem[20][11] ), .B2(n269), .ZN(
        n1445) );
  MAOI22D0 U1081 ( .A1(n269), .A2(n615), .B1(\mem[20][12] ), .B2(n269), .ZN(
        n1446) );
  MAOI22D0 U1082 ( .A1(n269), .A2(n373), .B1(\mem[20][13] ), .B2(n269), .ZN(
        n1447) );
  MAOI22D0 U1083 ( .A1(n269), .A2(n637), .B1(\mem[20][14] ), .B2(n269), .ZN(
        n1448) );
  MAOI22D0 U1084 ( .A1(n269), .A2(n351), .B1(\mem[20][15] ), .B2(n269), .ZN(
        n1449) );
  MAOI22D0 U1085 ( .A1(n269), .A2(n659), .B1(\mem[20][16] ), .B2(n269), .ZN(
        n1450) );
  MAOI22D0 U1086 ( .A1(n269), .A2(n329), .B1(\mem[20][17] ), .B2(n269), .ZN(
        n1451) );
  MAOI22D0 U1087 ( .A1(n269), .A2(n681), .B1(\mem[20][18] ), .B2(n269), .ZN(
        n1452) );
  MAOI22D0 U1088 ( .A1(n269), .A2(n307), .B1(\mem[20][19] ), .B2(n269), .ZN(
        n1453) );
  MAOI22D0 U1089 ( .A1(n269), .A2(n285), .B1(\mem[20][21] ), .B2(n269), .ZN(
        n1455) );
  MAOI22D0 U1090 ( .A1(n269), .A2(n725), .B1(\mem[20][22] ), .B2(n269), .ZN(
        n1456) );
  MAOI22D0 U1091 ( .A1(n269), .A2(n279), .B1(\mem[20][23] ), .B2(n269), .ZN(
        n1457) );
  NR2XD0 U1092 ( .A1(n270), .A2(n277), .ZN(n271) );
  MAOI22D0 U1093 ( .A1(n271), .A2(n281), .B1(\mem[19][0] ), .B2(n271), .ZN(
        n1458) );
  MAOI22D0 U1094 ( .A1(n271), .A2(n505), .B1(\mem[19][1] ), .B2(n271), .ZN(
        n1459) );
  MAOI22D0 U1095 ( .A1(n271), .A2(n755), .B1(\mem[19][2] ), .B2(n271), .ZN(
        n1460) );
  MAOI22D0 U1096 ( .A1(n271), .A2(n483), .B1(\mem[19][3] ), .B2(n271), .ZN(
        n1461) );
  MAOI22D0 U1097 ( .A1(n271), .A2(n527), .B1(\mem[19][4] ), .B2(n271), .ZN(
        n1462) );
  MAOI22D0 U1098 ( .A1(n271), .A2(n461), .B1(\mem[19][5] ), .B2(n271), .ZN(
        n1463) );
  MAOI22D0 U1099 ( .A1(n271), .A2(n549), .B1(\mem[19][6] ), .B2(n271), .ZN(
        n1464) );
  MAOI22D0 U1100 ( .A1(n271), .A2(n439), .B1(\mem[19][7] ), .B2(n271), .ZN(
        n1465) );
  MAOI22D0 U1101 ( .A1(n271), .A2(n571), .B1(\mem[19][8] ), .B2(n271), .ZN(
        n1466) );
  MAOI22D0 U1102 ( .A1(n271), .A2(n417), .B1(\mem[19][9] ), .B2(n271), .ZN(
        n1467) );
  MAOI22D0 U1103 ( .A1(n271), .A2(n593), .B1(\mem[19][10] ), .B2(n271), .ZN(
        n1468) );
  MAOI22D0 U1104 ( .A1(n271), .A2(n615), .B1(\mem[19][12] ), .B2(n271), .ZN(
        n1470) );
  MAOI22D0 U1105 ( .A1(n271), .A2(n373), .B1(\mem[19][13] ), .B2(n271), .ZN(
        n1471) );
  MAOI22D0 U1106 ( .A1(n271), .A2(n637), .B1(\mem[19][14] ), .B2(n271), .ZN(
        n1472) );
  MAOI22D0 U1107 ( .A1(n271), .A2(n351), .B1(\mem[19][15] ), .B2(n271), .ZN(
        n1473) );
  MAOI22D0 U1108 ( .A1(n271), .A2(n659), .B1(\mem[19][16] ), .B2(n271), .ZN(
        n1474) );
  MAOI22D0 U1109 ( .A1(n271), .A2(n329), .B1(\mem[19][17] ), .B2(n271), .ZN(
        n1475) );
  MAOI22D0 U1110 ( .A1(n271), .A2(n681), .B1(\mem[19][18] ), .B2(n271), .ZN(
        n1476) );
  MAOI22D0 U1111 ( .A1(n271), .A2(n307), .B1(\mem[19][19] ), .B2(n271), .ZN(
        n1477) );
  MAOI22D0 U1112 ( .A1(n271), .A2(n703), .B1(\mem[19][20] ), .B2(n271), .ZN(
        n1478) );
  MAOI22D0 U1113 ( .A1(n271), .A2(n285), .B1(\mem[19][21] ), .B2(n271), .ZN(
        n1479) );
  MAOI22D0 U1114 ( .A1(n271), .A2(n725), .B1(\mem[19][22] ), .B2(n271), .ZN(
        n1480) );
  MAOI22D0 U1115 ( .A1(n271), .A2(n279), .B1(\mem[19][23] ), .B2(n271), .ZN(
        n1481) );
  NR2XD0 U1116 ( .A1(n272), .A2(n277), .ZN(n274) );
  MAOI22D0 U1117 ( .A1(n274), .A2(n281), .B1(\mem[18][0] ), .B2(n274), .ZN(
        n1482) );
  MAOI22D0 U1118 ( .A1(n274), .A2(n505), .B1(\mem[18][1] ), .B2(n274), .ZN(
        n1483) );
  MAOI22D0 U1119 ( .A1(n274), .A2(n483), .B1(\mem[18][3] ), .B2(n274), .ZN(
        n1485) );
  MAOI22D0 U1120 ( .A1(n274), .A2(n527), .B1(\mem[18][4] ), .B2(n274), .ZN(
        n1486) );
  MAOI22D0 U1121 ( .A1(n274), .A2(n461), .B1(\mem[18][5] ), .B2(n274), .ZN(
        n1487) );
  MAOI22D0 U1122 ( .A1(n274), .A2(n549), .B1(\mem[18][6] ), .B2(n274), .ZN(
        n1488) );
  MAOI22D0 U1123 ( .A1(n274), .A2(n439), .B1(\mem[18][7] ), .B2(n274), .ZN(
        n1489) );
  MAOI22D0 U1124 ( .A1(n274), .A2(n571), .B1(\mem[18][8] ), .B2(n274), .ZN(
        n1490) );
  MAOI22D0 U1125 ( .A1(n274), .A2(n417), .B1(\mem[18][9] ), .B2(n274), .ZN(
        n1491) );
  MAOI22D0 U1126 ( .A1(n274), .A2(n593), .B1(\mem[18][10] ), .B2(n274), .ZN(
        n1492) );
  MAOI22D0 U1127 ( .A1(n274), .A2(n395), .B1(\mem[18][11] ), .B2(n274), .ZN(
        n1493) );
  MAOI22D0 U1128 ( .A1(n274), .A2(n615), .B1(\mem[18][12] ), .B2(n274), .ZN(
        n1494) );
  MAOI22D0 U1129 ( .A1(n274), .A2(n373), .B1(\mem[18][13] ), .B2(n274), .ZN(
        n1495) );
  MAOI22D0 U1130 ( .A1(n273), .A2(n549), .B1(\mem[21][6] ), .B2(n273), .ZN(
        n1416) );
  MAOI22D0 U1131 ( .A1(n274), .A2(n637), .B1(\mem[18][14] ), .B2(n274), .ZN(
        n1496) );
  MAOI22D0 U1132 ( .A1(n274), .A2(n351), .B1(\mem[18][15] ), .B2(n274), .ZN(
        n1497) );
  MAOI22D0 U1133 ( .A1(n274), .A2(n659), .B1(\mem[18][16] ), .B2(n274), .ZN(
        n1498) );
  MAOI22D0 U1134 ( .A1(n274), .A2(n681), .B1(\mem[18][18] ), .B2(n274), .ZN(
        n1500) );
  MAOI22D0 U1135 ( .A1(n274), .A2(n307), .B1(\mem[18][19] ), .B2(n274), .ZN(
        n1501) );
  MAOI22D0 U1136 ( .A1(n274), .A2(n703), .B1(\mem[18][20] ), .B2(n274), .ZN(
        n1502) );
  MAOI22D0 U1137 ( .A1(n274), .A2(n285), .B1(\mem[18][21] ), .B2(n274), .ZN(
        n1503) );
  MAOI22D0 U1138 ( .A1(n274), .A2(n725), .B1(\mem[18][22] ), .B2(n274), .ZN(
        n1504) );
  MAOI22D0 U1139 ( .A1(n274), .A2(n279), .B1(\mem[18][23] ), .B2(n274), .ZN(
        n1505) );
  NR2XD0 U1140 ( .A1(n275), .A2(n277), .ZN(n276) );
  MAOI22D0 U1141 ( .A1(n276), .A2(n281), .B1(\mem[17][0] ), .B2(n276), .ZN(
        n1506) );
  MAOI22D0 U1142 ( .A1(n276), .A2(n505), .B1(\mem[17][1] ), .B2(n276), .ZN(
        n1507) );
  MAOI22D0 U1143 ( .A1(n276), .A2(n755), .B1(\mem[17][2] ), .B2(n276), .ZN(
        n1508) );
  MAOI22D0 U1144 ( .A1(n276), .A2(n483), .B1(\mem[17][3] ), .B2(n276), .ZN(
        n1509) );
  MAOI22D0 U1145 ( .A1(n276), .A2(n527), .B1(\mem[17][4] ), .B2(n276), .ZN(
        n1510) );
  MAOI22D0 U1146 ( .A1(n276), .A2(n461), .B1(\mem[17][5] ), .B2(n276), .ZN(
        n1511) );
  MAOI22D0 U1147 ( .A1(n276), .A2(n549), .B1(\mem[17][6] ), .B2(n276), .ZN(
        n1512) );
  MAOI22D0 U1148 ( .A1(n276), .A2(n439), .B1(\mem[17][7] ), .B2(n276), .ZN(
        n1513) );
  MAOI22D0 U1149 ( .A1(n276), .A2(n417), .B1(\mem[17][9] ), .B2(n276), .ZN(
        n1515) );
  MAOI22D0 U1150 ( .A1(n276), .A2(n593), .B1(\mem[17][10] ), .B2(n276), .ZN(
        n1516) );
  MAOI22D0 U1151 ( .A1(n276), .A2(n395), .B1(\mem[17][11] ), .B2(n276), .ZN(
        n1517) );
  MAOI22D0 U1152 ( .A1(n276), .A2(n615), .B1(\mem[17][12] ), .B2(n276), .ZN(
        n1518) );
  MAOI22D0 U1153 ( .A1(n276), .A2(n373), .B1(\mem[17][13] ), .B2(n276), .ZN(
        n1519) );
  MAOI22D0 U1154 ( .A1(n276), .A2(n637), .B1(\mem[17][14] ), .B2(n276), .ZN(
        n1520) );
  MAOI22D0 U1155 ( .A1(n276), .A2(n351), .B1(\mem[17][15] ), .B2(n276), .ZN(
        n1521) );
  MAOI22D0 U1156 ( .A1(n276), .A2(n659), .B1(\mem[17][16] ), .B2(n276), .ZN(
        n1522) );
  MAOI22D0 U1157 ( .A1(n276), .A2(n329), .B1(\mem[17][17] ), .B2(n276), .ZN(
        n1523) );
  MAOI22D0 U1158 ( .A1(n276), .A2(n681), .B1(\mem[17][18] ), .B2(n276), .ZN(
        n1524) );
  MAOI22D0 U1159 ( .A1(n276), .A2(n307), .B1(\mem[17][19] ), .B2(n276), .ZN(
        n1525) );
  MAOI22D0 U1160 ( .A1(n276), .A2(n703), .B1(\mem[17][20] ), .B2(n276), .ZN(
        n1526) );
  MAOI22D0 U1161 ( .A1(n276), .A2(n285), .B1(\mem[17][21] ), .B2(n276), .ZN(
        n1527) );
  MAOI22D0 U1162 ( .A1(n276), .A2(n725), .B1(\mem[17][22] ), .B2(n276), .ZN(
        n1528) );
  NR2XD0 U1163 ( .A1(n278), .A2(n277), .ZN(n280) );
  MAOI22D0 U1164 ( .A1(n280), .A2(n281), .B1(\mem[16][0] ), .B2(n280), .ZN(
        n1530) );
  MAOI22D0 U1165 ( .A1(n280), .A2(n505), .B1(\mem[16][1] ), .B2(n280), .ZN(
        n1531) );
  MAOI22D0 U1166 ( .A1(n280), .A2(n755), .B1(\mem[16][2] ), .B2(n280), .ZN(
        n1532) );
  MAOI22D0 U1167 ( .A1(n280), .A2(n483), .B1(\mem[16][3] ), .B2(n280), .ZN(
        n1533) );
  MAOI22D0 U1168 ( .A1(n280), .A2(n527), .B1(\mem[16][4] ), .B2(n280), .ZN(
        n1534) );
  MAOI22D0 U1169 ( .A1(n280), .A2(n461), .B1(\mem[16][5] ), .B2(n280), .ZN(
        n1535) );
  MAOI22D0 U1170 ( .A1(n280), .A2(n549), .B1(\mem[16][6] ), .B2(n280), .ZN(
        n1536) );
  MAOI22D0 U1171 ( .A1(n280), .A2(n439), .B1(\mem[16][7] ), .B2(n280), .ZN(
        n1537) );
  MAOI22D0 U1172 ( .A1(n280), .A2(n571), .B1(\mem[16][8] ), .B2(n280), .ZN(
        n1538) );
  MAOI22D0 U1173 ( .A1(n280), .A2(n417), .B1(\mem[16][9] ), .B2(n280), .ZN(
        n1539) );
  MAOI22D0 U1174 ( .A1(n280), .A2(n593), .B1(\mem[16][10] ), .B2(n280), .ZN(
        n1540) );
  MAOI22D0 U1175 ( .A1(n280), .A2(n395), .B1(\mem[16][11] ), .B2(n280), .ZN(
        n1541) );
  MAOI22D0 U1176 ( .A1(n280), .A2(n615), .B1(\mem[16][12] ), .B2(n280), .ZN(
        n1542) );
  MAOI22D0 U1177 ( .A1(n280), .A2(n373), .B1(\mem[16][13] ), .B2(n280), .ZN(
        n1543) );
  MAOI22D0 U1178 ( .A1(n280), .A2(n351), .B1(\mem[16][15] ), .B2(n280), .ZN(
        n1545) );
  MAOI22D0 U1179 ( .A1(n280), .A2(n659), .B1(\mem[16][16] ), .B2(n280), .ZN(
        n1546) );
  MAOI22D0 U1180 ( .A1(n280), .A2(n329), .B1(\mem[16][17] ), .B2(n280), .ZN(
        n1547) );
  MAOI22D0 U1181 ( .A1(n280), .A2(n681), .B1(\mem[16][18] ), .B2(n280), .ZN(
        n1548) );
  MAOI22D0 U1182 ( .A1(n280), .A2(n307), .B1(\mem[16][19] ), .B2(n280), .ZN(
        n1549) );
  MAOI22D0 U1183 ( .A1(n280), .A2(n703), .B1(\mem[16][20] ), .B2(n280), .ZN(
        n1550) );
  MAOI22D0 U1184 ( .A1(n280), .A2(n285), .B1(\mem[16][21] ), .B2(n280), .ZN(
        n1551) );
  MAOI22D0 U1185 ( .A1(n280), .A2(n725), .B1(\mem[16][22] ), .B2(n280), .ZN(
        n1552) );
  MAOI22D0 U1186 ( .A1(n280), .A2(n279), .B1(\mem[16][23] ), .B2(n280), .ZN(
        n1553) );
  MAOI22D0 U1187 ( .A1(n282), .A2(n281), .B1(\mem[15][0] ), .B2(n282), .ZN(
        n1554) );
  MAOI22D0 U1188 ( .A1(n282), .A2(n505), .B1(\mem[15][1] ), .B2(n282), .ZN(
        n1555) );
  MAOI22D0 U1189 ( .A1(n282), .A2(n755), .B1(\mem[15][2] ), .B2(n282), .ZN(
        n1556) );
  MAOI22D0 U1190 ( .A1(n282), .A2(n483), .B1(\mem[15][3] ), .B2(n282), .ZN(
        n1557) );
  MAOI22D0 U1191 ( .A1(n282), .A2(n527), .B1(\mem[15][4] ), .B2(n282), .ZN(
        n1558) );
  MAOI22D0 U1192 ( .A1(n282), .A2(n549), .B1(\mem[15][6] ), .B2(n282), .ZN(
        n1560) );
  MAOI22D0 U1193 ( .A1(n282), .A2(n439), .B1(\mem[15][7] ), .B2(n282), .ZN(
        n1561) );
  MAOI22D0 U1194 ( .A1(n282), .A2(n571), .B1(\mem[15][8] ), .B2(n282), .ZN(
        n1562) );
  MAOI22D0 U1195 ( .A1(n282), .A2(n417), .B1(\mem[15][9] ), .B2(n282), .ZN(
        n1563) );
  MAOI22D0 U1196 ( .A1(n282), .A2(n593), .B1(\mem[15][10] ), .B2(n282), .ZN(
        n1564) );
  MAOI22D0 U1197 ( .A1(n282), .A2(n395), .B1(\mem[15][11] ), .B2(n282), .ZN(
        n1565) );
  MAOI22D0 U1198 ( .A1(n282), .A2(n615), .B1(\mem[15][12] ), .B2(n282), .ZN(
        n1566) );
  MAOI22D0 U1199 ( .A1(n282), .A2(n373), .B1(\mem[15][13] ), .B2(n282), .ZN(
        n1567) );
  MAOI22D0 U1200 ( .A1(n282), .A2(n637), .B1(\mem[15][14] ), .B2(n282), .ZN(
        n1568) );
  MAOI22D0 U1201 ( .A1(n282), .A2(n351), .B1(\mem[15][15] ), .B2(n282), .ZN(
        n1569) );
  MAOI22D0 U1202 ( .A1(n282), .A2(n659), .B1(\mem[15][16] ), .B2(n282), .ZN(
        n1570) );
  MAOI22D0 U1203 ( .A1(n282), .A2(n329), .B1(\mem[15][17] ), .B2(n282), .ZN(
        n1571) );
  MAOI22D0 U1204 ( .A1(n282), .A2(n681), .B1(\mem[15][18] ), .B2(n282), .ZN(
        n1572) );
  AOI22D0 U1205 ( .A1(n746), .A2(\mem[30][21] ), .B1(n745), .B2(\mem[2][21] ), 
        .ZN(n304) );
  AOI22D0 U1206 ( .A1(n750), .A2(\mem[8][21] ), .B1(n749), .B2(\mem[10][21] ), 
        .ZN(n284) );
  AOI22D0 U1207 ( .A1(n752), .A2(\mem[6][21] ), .B1(n751), .B2(\mem[9][21] ), 
        .ZN(n283) );
  OA211D0 U1208 ( .A1(n756), .A2(n285), .B(n284), .C(n283), .Z(n302) );
  AOI22D0 U1209 ( .A1(n758), .A2(\mem[11][21] ), .B1(n757), .B2(\mem[4][21] ), 
        .ZN(n289) );
  AOI22D0 U1210 ( .A1(n760), .A2(\mem[5][21] ), .B1(n759), .B2(\mem[7][21] ), 
        .ZN(n288) );
  AOI22D0 U1211 ( .A1(n762), .A2(\mem[12][21] ), .B1(n761), .B2(\mem[14][21] ), 
        .ZN(n287) );
  AOI22D0 U1212 ( .A1(n764), .A2(\mem[13][21] ), .B1(n763), .B2(\mem[15][21] ), 
        .ZN(n286) );
  ND4D0 U1213 ( .A1(n289), .A2(n288), .A3(n287), .A4(n286), .ZN(n300) );
  AOI22D0 U1214 ( .A1(n770), .A2(\mem[16][21] ), .B1(n769), .B2(\mem[18][21] ), 
        .ZN(n293) );
  AOI22D0 U1215 ( .A1(n772), .A2(\mem[17][21] ), .B1(n771), .B2(\mem[19][21] ), 
        .ZN(n292) );
  AOI22D0 U1216 ( .A1(n776), .A2(\mem[25][21] ), .B1(n775), .B2(\mem[27][21] ), 
        .ZN(n290) );
  ND4D0 U1217 ( .A1(n293), .A2(n292), .A3(n291), .A4(n290), .ZN(n299) );
  AOI22D0 U1218 ( .A1(n782), .A2(\mem[20][21] ), .B1(n781), .B2(\mem[22][21] ), 
        .ZN(n297) );
  AOI22D0 U1219 ( .A1(n784), .A2(\mem[21][21] ), .B1(n783), .B2(\mem[23][21] ), 
        .ZN(n296) );
  AOI22D0 U1220 ( .A1(n786), .A2(\mem[28][21] ), .B1(n785), .B2(\mem[29][21] ), 
        .ZN(n295) );
  AOI22D0 U1221 ( .A1(n788), .A2(\mem[31][21] ), .B1(n787), .B2(\mem[0][21] ), 
        .ZN(n294) );
  NR3D0 U1222 ( .A1(n300), .A2(n299), .A3(n298), .ZN(n301) );
  ND4D0 U1223 ( .A1(n304), .A2(n303), .A3(n302), .A4(n301), .ZN(B[21]) );
  AOI22D0 U1224 ( .A1(n746), .A2(\mem[30][19] ), .B1(n745), .B2(\mem[2][19] ), 
        .ZN(n326) );
  AOI22D0 U1225 ( .A1(n748), .A2(\mem[1][19] ), .B1(n747), .B2(\mem[3][19] ), 
        .ZN(n325) );
  AOI22D0 U1226 ( .A1(n750), .A2(\mem[8][19] ), .B1(n749), .B2(\mem[10][19] ), 
        .ZN(n306) );
  AOI22D0 U1227 ( .A1(n752), .A2(\mem[6][19] ), .B1(n751), .B2(\mem[9][19] ), 
        .ZN(n305) );
  OA211D0 U1228 ( .A1(n756), .A2(n307), .B(n306), .C(n305), .Z(n324) );
  AOI22D0 U1229 ( .A1(n758), .A2(\mem[11][19] ), .B1(n757), .B2(\mem[4][19] ), 
        .ZN(n311) );
  AOI22D0 U1230 ( .A1(n760), .A2(\mem[5][19] ), .B1(n759), .B2(\mem[7][19] ), 
        .ZN(n310) );
  AOI22D0 U1231 ( .A1(n762), .A2(\mem[12][19] ), .B1(n761), .B2(\mem[14][19] ), 
        .ZN(n309) );
  AOI22D0 U1232 ( .A1(n764), .A2(\mem[13][19] ), .B1(n763), .B2(\mem[15][19] ), 
        .ZN(n308) );
  ND4D0 U1233 ( .A1(n311), .A2(n310), .A3(n309), .A4(n308), .ZN(n322) );
  AOI22D0 U1234 ( .A1(n770), .A2(\mem[16][19] ), .B1(n769), .B2(\mem[18][19] ), 
        .ZN(n315) );
  AOI22D0 U1235 ( .A1(n772), .A2(\mem[17][19] ), .B1(n771), .B2(\mem[19][19] ), 
        .ZN(n314) );
  AOI22D0 U1236 ( .A1(n774), .A2(\mem[24][19] ), .B1(n773), .B2(\mem[26][19] ), 
        .ZN(n313) );
  AOI22D0 U1237 ( .A1(n776), .A2(\mem[25][19] ), .B1(n775), .B2(\mem[27][19] ), 
        .ZN(n312) );
  ND4D0 U1238 ( .A1(n315), .A2(n314), .A3(n313), .A4(n312), .ZN(n321) );
  AOI22D0 U1239 ( .A1(n782), .A2(\mem[20][19] ), .B1(n781), .B2(\mem[22][19] ), 
        .ZN(n319) );
  AOI22D0 U1240 ( .A1(n784), .A2(\mem[21][19] ), .B1(n783), .B2(\mem[23][19] ), 
        .ZN(n318) );
  AOI22D0 U1241 ( .A1(n786), .A2(\mem[28][19] ), .B1(n785), .B2(\mem[29][19] ), 
        .ZN(n317) );
  AOI22D0 U1242 ( .A1(n788), .A2(\mem[31][19] ), .B1(n787), .B2(\mem[0][19] ), 
        .ZN(n316) );
  ND4D0 U1243 ( .A1(n319), .A2(n318), .A3(n317), .A4(n316), .ZN(n320) );
  NR3D0 U1244 ( .A1(n322), .A2(n321), .A3(n320), .ZN(n323) );
  ND4D0 U1245 ( .A1(n326), .A2(n325), .A3(n324), .A4(n323), .ZN(B[19]) );
  AOI22D0 U1246 ( .A1(n748), .A2(\mem[1][17] ), .B1(n747), .B2(\mem[3][17] ), 
        .ZN(n347) );
  AOI22D0 U1247 ( .A1(n750), .A2(\mem[8][17] ), .B1(n749), .B2(\mem[10][17] ), 
        .ZN(n328) );
  AOI22D0 U1248 ( .A1(n752), .A2(\mem[6][17] ), .B1(n751), .B2(\mem[9][17] ), 
        .ZN(n327) );
  OA211D0 U1249 ( .A1(n756), .A2(n329), .B(n328), .C(n327), .Z(n346) );
  AOI22D0 U1250 ( .A1(n758), .A2(\mem[11][17] ), .B1(n757), .B2(\mem[4][17] ), 
        .ZN(n333) );
  AOI22D0 U1251 ( .A1(n760), .A2(\mem[5][17] ), .B1(n759), .B2(\mem[7][17] ), 
        .ZN(n332) );
  AOI22D0 U1252 ( .A1(n762), .A2(\mem[12][17] ), .B1(n761), .B2(\mem[14][17] ), 
        .ZN(n331) );
  ND4D0 U1253 ( .A1(n333), .A2(n332), .A3(n331), .A4(n330), .ZN(n344) );
  AOI22D0 U1254 ( .A1(n770), .A2(\mem[16][17] ), .B1(n769), .B2(\mem[18][17] ), 
        .ZN(n337) );
  AOI22D0 U1255 ( .A1(n772), .A2(\mem[17][17] ), .B1(n771), .B2(\mem[19][17] ), 
        .ZN(n336) );
  AOI22D0 U1256 ( .A1(n774), .A2(\mem[24][17] ), .B1(n773), .B2(\mem[26][17] ), 
        .ZN(n335) );
  AOI22D0 U1257 ( .A1(n776), .A2(\mem[25][17] ), .B1(n775), .B2(\mem[27][17] ), 
        .ZN(n334) );
  ND4D0 U1258 ( .A1(n337), .A2(n336), .A3(n335), .A4(n334), .ZN(n343) );
  AOI22D0 U1259 ( .A1(n782), .A2(\mem[20][17] ), .B1(n781), .B2(\mem[22][17] ), 
        .ZN(n341) );
  AOI22D0 U1260 ( .A1(n784), .A2(\mem[21][17] ), .B1(n783), .B2(\mem[23][17] ), 
        .ZN(n340) );
  AOI22D0 U1261 ( .A1(n786), .A2(\mem[28][17] ), .B1(n785), .B2(\mem[29][17] ), 
        .ZN(n339) );
  AOI22D0 U1262 ( .A1(n788), .A2(\mem[31][17] ), .B1(n787), .B2(\mem[0][17] ), 
        .ZN(n338) );
  ND4D0 U1263 ( .A1(n341), .A2(n340), .A3(n339), .A4(n338), .ZN(n342) );
  NR3D0 U1264 ( .A1(n344), .A2(n343), .A3(n342), .ZN(n345) );
  ND4D0 U1265 ( .A1(n348), .A2(n347), .A3(n346), .A4(n345), .ZN(B[17]) );
  AOI22D0 U1266 ( .A1(n746), .A2(\mem[30][15] ), .B1(n745), .B2(\mem[2][15] ), 
        .ZN(n370) );
  AOI22D0 U1267 ( .A1(n748), .A2(\mem[1][15] ), .B1(n747), .B2(\mem[3][15] ), 
        .ZN(n369) );
  AOI22D0 U1268 ( .A1(n750), .A2(\mem[8][15] ), .B1(n749), .B2(\mem[10][15] ), 
        .ZN(n350) );
  AOI22D0 U1269 ( .A1(n752), .A2(\mem[6][15] ), .B1(n751), .B2(\mem[9][15] ), 
        .ZN(n349) );
  OA211D0 U1270 ( .A1(n756), .A2(n351), .B(n350), .C(n349), .Z(n368) );
  AOI22D0 U1271 ( .A1(n758), .A2(\mem[11][15] ), .B1(n757), .B2(\mem[4][15] ), 
        .ZN(n355) );
  AOI22D0 U1272 ( .A1(n760), .A2(\mem[5][15] ), .B1(n759), .B2(\mem[7][15] ), 
        .ZN(n354) );
  AOI22D0 U1273 ( .A1(n762), .A2(\mem[12][15] ), .B1(n761), .B2(\mem[14][15] ), 
        .ZN(n353) );
  AOI22D0 U1274 ( .A1(n764), .A2(\mem[13][15] ), .B1(n763), .B2(\mem[15][15] ), 
        .ZN(n352) );
  ND4D0 U1275 ( .A1(n355), .A2(n354), .A3(n353), .A4(n352), .ZN(n366) );
  AOI22D0 U1276 ( .A1(n770), .A2(\mem[16][15] ), .B1(n769), .B2(\mem[18][15] ), 
        .ZN(n359) );
  AOI22D0 U1277 ( .A1(n772), .A2(\mem[17][15] ), .B1(n771), .B2(\mem[19][15] ), 
        .ZN(n358) );
  AOI22D0 U1278 ( .A1(n774), .A2(\mem[24][15] ), .B1(n773), .B2(\mem[26][15] ), 
        .ZN(n357) );
  AOI22D0 U1279 ( .A1(n776), .A2(\mem[25][15] ), .B1(n775), .B2(\mem[27][15] ), 
        .ZN(n356) );
  ND4D0 U1280 ( .A1(n359), .A2(n358), .A3(n357), .A4(n356), .ZN(n365) );
  AOI22D0 U1281 ( .A1(n782), .A2(\mem[20][15] ), .B1(n781), .B2(\mem[22][15] ), 
        .ZN(n363) );
  AOI22D0 U1282 ( .A1(n786), .A2(\mem[28][15] ), .B1(n785), .B2(\mem[29][15] ), 
        .ZN(n361) );
  AOI22D0 U1283 ( .A1(n788), .A2(\mem[31][15] ), .B1(n787), .B2(\mem[0][15] ), 
        .ZN(n360) );
  NR3D0 U1284 ( .A1(n366), .A2(n365), .A3(n364), .ZN(n367) );
  ND4D0 U1285 ( .A1(n370), .A2(n369), .A3(n368), .A4(n367), .ZN(B[15]) );
  AOI22D0 U1286 ( .A1(n746), .A2(\mem[30][13] ), .B1(n745), .B2(\mem[2][13] ), 
        .ZN(n392) );
  AOI22D0 U1287 ( .A1(n748), .A2(\mem[1][13] ), .B1(n747), .B2(\mem[3][13] ), 
        .ZN(n391) );
  AOI22D0 U1288 ( .A1(n750), .A2(\mem[8][13] ), .B1(n749), .B2(\mem[10][13] ), 
        .ZN(n372) );
  AOI22D0 U1289 ( .A1(n752), .A2(\mem[6][13] ), .B1(n751), .B2(\mem[9][13] ), 
        .ZN(n371) );
  OA211D0 U1290 ( .A1(n756), .A2(n373), .B(n372), .C(n371), .Z(n390) );
  AOI22D0 U1291 ( .A1(n760), .A2(\mem[5][13] ), .B1(n759), .B2(\mem[7][13] ), 
        .ZN(n376) );
  AOI22D0 U1292 ( .A1(n762), .A2(\mem[12][13] ), .B1(n761), .B2(\mem[14][13] ), 
        .ZN(n375) );
  AOI22D0 U1293 ( .A1(n764), .A2(\mem[13][13] ), .B1(n763), .B2(\mem[15][13] ), 
        .ZN(n374) );
  ND4D0 U1294 ( .A1(n377), .A2(n376), .A3(n375), .A4(n374), .ZN(n388) );
  AOI22D0 U1295 ( .A1(n770), .A2(\mem[16][13] ), .B1(n769), .B2(\mem[18][13] ), 
        .ZN(n381) );
  AOI22D0 U1296 ( .A1(n772), .A2(\mem[17][13] ), .B1(n771), .B2(\mem[19][13] ), 
        .ZN(n380) );
  AOI22D0 U1297 ( .A1(n774), .A2(\mem[24][13] ), .B1(n773), .B2(\mem[26][13] ), 
        .ZN(n379) );
  AOI22D0 U1298 ( .A1(n776), .A2(\mem[25][13] ), .B1(n775), .B2(\mem[27][13] ), 
        .ZN(n378) );
  ND4D0 U1299 ( .A1(n381), .A2(n380), .A3(n379), .A4(n378), .ZN(n387) );
  AOI22D0 U1300 ( .A1(n782), .A2(\mem[20][13] ), .B1(n781), .B2(\mem[22][13] ), 
        .ZN(n385) );
  AOI22D0 U1301 ( .A1(n784), .A2(\mem[21][13] ), .B1(n783), .B2(\mem[23][13] ), 
        .ZN(n384) );
  AOI22D0 U1302 ( .A1(n786), .A2(\mem[28][13] ), .B1(n785), .B2(\mem[29][13] ), 
        .ZN(n383) );
  AOI22D0 U1303 ( .A1(n788), .A2(\mem[31][13] ), .B1(n787), .B2(\mem[0][13] ), 
        .ZN(n382) );
  ND4D0 U1304 ( .A1(n385), .A2(n384), .A3(n383), .A4(n382), .ZN(n386) );
  NR3D0 U1305 ( .A1(n388), .A2(n387), .A3(n386), .ZN(n389) );
  ND4D0 U1306 ( .A1(n392), .A2(n391), .A3(n390), .A4(n389), .ZN(B[13]) );
  AOI22D0 U1307 ( .A1(n746), .A2(\mem[30][11] ), .B1(n745), .B2(\mem[2][11] ), 
        .ZN(n414) );
  AOI22D0 U1308 ( .A1(n748), .A2(\mem[1][11] ), .B1(n747), .B2(\mem[3][11] ), 
        .ZN(n413) );
  AOI22D0 U1309 ( .A1(n750), .A2(\mem[8][11] ), .B1(n749), .B2(\mem[10][11] ), 
        .ZN(n394) );
  AOI22D0 U1310 ( .A1(n752), .A2(\mem[6][11] ), .B1(n751), .B2(\mem[9][11] ), 
        .ZN(n393) );
  OA211D0 U1311 ( .A1(n756), .A2(n395), .B(n394), .C(n393), .Z(n412) );
  AOI22D0 U1312 ( .A1(n758), .A2(\mem[11][11] ), .B1(n757), .B2(\mem[4][11] ), 
        .ZN(n399) );
  AOI22D0 U1313 ( .A1(n760), .A2(\mem[5][11] ), .B1(n759), .B2(\mem[7][11] ), 
        .ZN(n398) );
  AOI22D0 U1314 ( .A1(n762), .A2(\mem[12][11] ), .B1(n761), .B2(\mem[14][11] ), 
        .ZN(n397) );
  AOI22D0 U1315 ( .A1(n764), .A2(\mem[13][11] ), .B1(n763), .B2(\mem[15][11] ), 
        .ZN(n396) );
  ND4D0 U1316 ( .A1(n399), .A2(n398), .A3(n397), .A4(n396), .ZN(n410) );
  AOI22D0 U1317 ( .A1(n770), .A2(\mem[16][11] ), .B1(n769), .B2(\mem[18][11] ), 
        .ZN(n403) );
  AOI22D0 U1318 ( .A1(n772), .A2(\mem[17][11] ), .B1(n771), .B2(\mem[19][11] ), 
        .ZN(n402) );
  AOI22D0 U1319 ( .A1(n776), .A2(\mem[25][11] ), .B1(n775), .B2(\mem[27][11] ), 
        .ZN(n400) );
  ND4D0 U1320 ( .A1(n403), .A2(n402), .A3(n401), .A4(n400), .ZN(n409) );
  AOI22D0 U1321 ( .A1(n782), .A2(\mem[20][11] ), .B1(n781), .B2(\mem[22][11] ), 
        .ZN(n407) );
  AOI22D0 U1322 ( .A1(n784), .A2(\mem[21][11] ), .B1(n783), .B2(\mem[23][11] ), 
        .ZN(n406) );
  AOI22D0 U1323 ( .A1(n786), .A2(\mem[28][11] ), .B1(n785), .B2(\mem[29][11] ), 
        .ZN(n405) );
  AOI22D0 U1324 ( .A1(n788), .A2(\mem[31][11] ), .B1(n787), .B2(\mem[0][11] ), 
        .ZN(n404) );
  ND4D0 U1325 ( .A1(n407), .A2(n406), .A3(n405), .A4(n404), .ZN(n408) );
  NR3D0 U1326 ( .A1(n410), .A2(n409), .A3(n408), .ZN(n411) );
  ND4D0 U1327 ( .A1(n414), .A2(n413), .A3(n412), .A4(n411), .ZN(B[11]) );
  AOI22D0 U1328 ( .A1(n746), .A2(\mem[30][9] ), .B1(n745), .B2(\mem[2][9] ), 
        .ZN(n436) );
  AOI22D0 U1329 ( .A1(n748), .A2(\mem[1][9] ), .B1(n747), .B2(\mem[3][9] ), 
        .ZN(n435) );
  AOI22D0 U1330 ( .A1(n750), .A2(\mem[8][9] ), .B1(n749), .B2(\mem[10][9] ), 
        .ZN(n416) );
  AOI22D0 U1331 ( .A1(n752), .A2(\mem[6][9] ), .B1(n751), .B2(\mem[9][9] ), 
        .ZN(n415) );
  OA211D0 U1332 ( .A1(n756), .A2(n417), .B(n416), .C(n415), .Z(n434) );
  AOI22D0 U1333 ( .A1(n758), .A2(\mem[11][9] ), .B1(n757), .B2(\mem[4][9] ), 
        .ZN(n421) );
  AOI22D0 U1334 ( .A1(n760), .A2(\mem[5][9] ), .B1(n759), .B2(\mem[7][9] ), 
        .ZN(n420) );
  AOI22D0 U1335 ( .A1(n762), .A2(\mem[12][9] ), .B1(n761), .B2(\mem[14][9] ), 
        .ZN(n419) );
  AOI22D0 U1336 ( .A1(n764), .A2(\mem[13][9] ), .B1(n763), .B2(\mem[15][9] ), 
        .ZN(n418) );
  ND4D0 U1337 ( .A1(n421), .A2(n420), .A3(n419), .A4(n418), .ZN(n432) );
  AOI22D0 U1338 ( .A1(n770), .A2(\mem[16][9] ), .B1(n769), .B2(\mem[18][9] ), 
        .ZN(n425) );
  AOI22D0 U1339 ( .A1(n772), .A2(\mem[17][9] ), .B1(n771), .B2(\mem[19][9] ), 
        .ZN(n424) );
  AOI22D0 U1340 ( .A1(n774), .A2(\mem[24][9] ), .B1(n773), .B2(\mem[26][9] ), 
        .ZN(n423) );
  AOI22D0 U1341 ( .A1(n776), .A2(\mem[25][9] ), .B1(n775), .B2(\mem[27][9] ), 
        .ZN(n422) );
  ND4D0 U1342 ( .A1(n425), .A2(n424), .A3(n423), .A4(n422), .ZN(n431) );
  AOI22D0 U1343 ( .A1(n782), .A2(\mem[20][9] ), .B1(n781), .B2(\mem[22][9] ), 
        .ZN(n429) );
  AOI22D0 U1344 ( .A1(n784), .A2(\mem[21][9] ), .B1(n783), .B2(\mem[23][9] ), 
        .ZN(n428) );
  AOI22D0 U1345 ( .A1(n786), .A2(\mem[28][9] ), .B1(n785), .B2(\mem[29][9] ), 
        .ZN(n427) );
  AOI22D0 U1346 ( .A1(n788), .A2(\mem[31][9] ), .B1(n787), .B2(\mem[0][9] ), 
        .ZN(n426) );
  NR3D0 U1347 ( .A1(n432), .A2(n431), .A3(n430), .ZN(n433) );
  ND4D0 U1348 ( .A1(n436), .A2(n435), .A3(n434), .A4(n433), .ZN(B[9]) );
  AOI22D0 U1349 ( .A1(n746), .A2(\mem[30][7] ), .B1(n745), .B2(\mem[2][7] ), 
        .ZN(n458) );
  AOI22D0 U1350 ( .A1(n748), .A2(\mem[1][7] ), .B1(n747), .B2(\mem[3][7] ), 
        .ZN(n457) );
  AOI22D0 U1351 ( .A1(n750), .A2(\mem[8][7] ), .B1(n749), .B2(\mem[10][7] ), 
        .ZN(n438) );
  AOI22D0 U1352 ( .A1(n752), .A2(\mem[6][7] ), .B1(n751), .B2(\mem[9][7] ), 
        .ZN(n437) );
  OA211D0 U1353 ( .A1(n756), .A2(n439), .B(n438), .C(n437), .Z(n456) );
  AOI22D0 U1354 ( .A1(n758), .A2(\mem[11][7] ), .B1(n757), .B2(\mem[4][7] ), 
        .ZN(n443) );
  AOI22D0 U1355 ( .A1(n760), .A2(\mem[5][7] ), .B1(n759), .B2(\mem[7][7] ), 
        .ZN(n442) );
  AOI22D0 U1356 ( .A1(n762), .A2(\mem[12][7] ), .B1(n761), .B2(\mem[14][7] ), 
        .ZN(n441) );
  ND4D0 U1357 ( .A1(n443), .A2(n442), .A3(n441), .A4(n440), .ZN(n454) );
  AOI22D0 U1358 ( .A1(n770), .A2(\mem[16][7] ), .B1(n769), .B2(\mem[18][7] ), 
        .ZN(n447) );
  AOI22D0 U1359 ( .A1(n772), .A2(\mem[17][7] ), .B1(n771), .B2(\mem[19][7] ), 
        .ZN(n446) );
  AOI22D0 U1360 ( .A1(n774), .A2(\mem[24][7] ), .B1(n773), .B2(\mem[26][7] ), 
        .ZN(n445) );
  AOI22D0 U1361 ( .A1(n776), .A2(\mem[25][7] ), .B1(n775), .B2(\mem[27][7] ), 
        .ZN(n444) );
  ND4D0 U1362 ( .A1(n447), .A2(n446), .A3(n445), .A4(n444), .ZN(n453) );
  AOI22D0 U1363 ( .A1(n782), .A2(\mem[20][7] ), .B1(n781), .B2(\mem[22][7] ), 
        .ZN(n451) );
  AOI22D0 U1364 ( .A1(n784), .A2(\mem[21][7] ), .B1(n783), .B2(\mem[23][7] ), 
        .ZN(n450) );
  AOI22D0 U1365 ( .A1(n786), .A2(\mem[28][7] ), .B1(n785), .B2(\mem[29][7] ), 
        .ZN(n449) );
  AOI22D0 U1366 ( .A1(n788), .A2(\mem[31][7] ), .B1(n787), .B2(\mem[0][7] ), 
        .ZN(n448) );
  ND4D0 U1367 ( .A1(n451), .A2(n450), .A3(n449), .A4(n448), .ZN(n452) );
  NR3D0 U1368 ( .A1(n454), .A2(n453), .A3(n452), .ZN(n455) );
  AOI22D0 U1369 ( .A1(n746), .A2(\mem[30][5] ), .B1(n745), .B2(\mem[2][5] ), 
        .ZN(n480) );
  AOI22D0 U1370 ( .A1(n748), .A2(\mem[1][5] ), .B1(n747), .B2(\mem[3][5] ), 
        .ZN(n479) );
  AOI22D0 U1371 ( .A1(n750), .A2(\mem[8][5] ), .B1(n749), .B2(\mem[10][5] ), 
        .ZN(n460) );
  AOI22D0 U1372 ( .A1(n752), .A2(\mem[6][5] ), .B1(n751), .B2(\mem[9][5] ), 
        .ZN(n459) );
  OA211D0 U1373 ( .A1(n756), .A2(n461), .B(n460), .C(n459), .Z(n478) );
  AOI22D0 U1374 ( .A1(n758), .A2(\mem[11][5] ), .B1(n757), .B2(\mem[4][5] ), 
        .ZN(n465) );
  AOI22D0 U1375 ( .A1(n760), .A2(\mem[5][5] ), .B1(n759), .B2(\mem[7][5] ), 
        .ZN(n464) );
  AOI22D0 U1376 ( .A1(n762), .A2(\mem[12][5] ), .B1(n761), .B2(\mem[14][5] ), 
        .ZN(n463) );
  AOI22D0 U1377 ( .A1(n764), .A2(\mem[13][5] ), .B1(n763), .B2(\mem[15][5] ), 
        .ZN(n462) );
  ND4D0 U1378 ( .A1(n465), .A2(n464), .A3(n463), .A4(n462), .ZN(n476) );
  AOI22D0 U1379 ( .A1(n770), .A2(\mem[16][5] ), .B1(n769), .B2(\mem[18][5] ), 
        .ZN(n469) );
  AOI22D0 U1380 ( .A1(n772), .A2(\mem[17][5] ), .B1(n771), .B2(\mem[19][5] ), 
        .ZN(n468) );
  AOI22D0 U1381 ( .A1(n774), .A2(\mem[24][5] ), .B1(n773), .B2(\mem[26][5] ), 
        .ZN(n467) );
  AOI22D0 U1382 ( .A1(n776), .A2(\mem[25][5] ), .B1(n775), .B2(\mem[27][5] ), 
        .ZN(n466) );
  ND4D0 U1383 ( .A1(n469), .A2(n468), .A3(n467), .A4(n466), .ZN(n475) );
  AOI22D0 U1384 ( .A1(n782), .A2(\mem[20][5] ), .B1(n781), .B2(\mem[22][5] ), 
        .ZN(n473) );
  AOI22D0 U1385 ( .A1(n786), .A2(\mem[28][5] ), .B1(n785), .B2(\mem[29][5] ), 
        .ZN(n471) );
  AOI22D0 U1386 ( .A1(n788), .A2(\mem[31][5] ), .B1(n787), .B2(\mem[0][5] ), 
        .ZN(n470) );
  ND4D0 U1387 ( .A1(n473), .A2(n472), .A3(n471), .A4(n470), .ZN(n474) );
  NR3D0 U1388 ( .A1(n476), .A2(n475), .A3(n474), .ZN(n477) );
  ND4D0 U1389 ( .A1(n480), .A2(n479), .A3(n478), .A4(n477), .ZN(B[5]) );
  AOI22D0 U1390 ( .A1(n746), .A2(\mem[30][3] ), .B1(n745), .B2(\mem[2][3] ), 
        .ZN(n502) );
  AOI22D0 U1391 ( .A1(n748), .A2(\mem[1][3] ), .B1(n747), .B2(\mem[3][3] ), 
        .ZN(n501) );
  AOI22D0 U1392 ( .A1(n750), .A2(\mem[8][3] ), .B1(n749), .B2(\mem[10][3] ), 
        .ZN(n482) );
  AOI22D0 U1393 ( .A1(n752), .A2(\mem[6][3] ), .B1(n751), .B2(\mem[9][3] ), 
        .ZN(n481) );
  OA211D0 U1394 ( .A1(n756), .A2(n483), .B(n482), .C(n481), .Z(n500) );
  AOI22D0 U1395 ( .A1(n760), .A2(\mem[5][3] ), .B1(n759), .B2(\mem[7][3] ), 
        .ZN(n486) );
  AOI22D0 U1396 ( .A1(n762), .A2(\mem[12][3] ), .B1(n761), .B2(\mem[14][3] ), 
        .ZN(n485) );
  AOI22D0 U1397 ( .A1(n764), .A2(\mem[13][3] ), .B1(n763), .B2(\mem[15][3] ), 
        .ZN(n484) );
  ND4D0 U1398 ( .A1(n487), .A2(n486), .A3(n485), .A4(n484), .ZN(n498) );
  AOI22D0 U1399 ( .A1(n770), .A2(\mem[16][3] ), .B1(n769), .B2(\mem[18][3] ), 
        .ZN(n491) );
  AOI22D0 U1400 ( .A1(n772), .A2(\mem[17][3] ), .B1(n771), .B2(\mem[19][3] ), 
        .ZN(n490) );
  AOI22D0 U1401 ( .A1(n774), .A2(\mem[24][3] ), .B1(n773), .B2(\mem[26][3] ), 
        .ZN(n489) );
  AOI22D0 U1402 ( .A1(n776), .A2(\mem[25][3] ), .B1(n775), .B2(\mem[27][3] ), 
        .ZN(n488) );
  ND4D0 U1403 ( .A1(n491), .A2(n490), .A3(n489), .A4(n488), .ZN(n497) );
  AOI22D0 U1404 ( .A1(n782), .A2(\mem[20][3] ), .B1(n781), .B2(\mem[22][3] ), 
        .ZN(n495) );
  AOI22D0 U1405 ( .A1(n784), .A2(\mem[21][3] ), .B1(n783), .B2(\mem[23][3] ), 
        .ZN(n494) );
  AOI22D0 U1406 ( .A1(n786), .A2(\mem[28][3] ), .B1(n785), .B2(\mem[29][3] ), 
        .ZN(n493) );
  AOI22D0 U1407 ( .A1(n788), .A2(\mem[31][3] ), .B1(n787), .B2(\mem[0][3] ), 
        .ZN(n492) );
  NR3D0 U1408 ( .A1(n498), .A2(n497), .A3(n496), .ZN(n499) );
  ND4D0 U1409 ( .A1(n502), .A2(n501), .A3(n500), .A4(n499), .ZN(B[3]) );
  AOI22D0 U1410 ( .A1(n746), .A2(\mem[30][1] ), .B1(n745), .B2(\mem[2][1] ), 
        .ZN(n524) );
  AOI22D0 U1411 ( .A1(n748), .A2(\mem[1][1] ), .B1(n747), .B2(\mem[3][1] ), 
        .ZN(n523) );
  AOI22D0 U1412 ( .A1(n750), .A2(\mem[8][1] ), .B1(n749), .B2(\mem[10][1] ), 
        .ZN(n504) );
  AOI22D0 U1413 ( .A1(n752), .A2(\mem[6][1] ), .B1(n751), .B2(\mem[9][1] ), 
        .ZN(n503) );
  OA211D0 U1414 ( .A1(n756), .A2(n505), .B(n504), .C(n503), .Z(n522) );
  AOI22D0 U1415 ( .A1(n758), .A2(\mem[11][1] ), .B1(n757), .B2(\mem[4][1] ), 
        .ZN(n509) );
  AOI22D0 U1416 ( .A1(n760), .A2(\mem[5][1] ), .B1(n759), .B2(\mem[7][1] ), 
        .ZN(n508) );
  AOI22D0 U1417 ( .A1(n762), .A2(\mem[12][1] ), .B1(n761), .B2(\mem[14][1] ), 
        .ZN(n507) );
  AOI22D0 U1418 ( .A1(n764), .A2(\mem[13][1] ), .B1(n763), .B2(\mem[15][1] ), 
        .ZN(n506) );
  ND4D0 U1419 ( .A1(n509), .A2(n508), .A3(n507), .A4(n506), .ZN(n520) );
  AOI22D0 U1420 ( .A1(n770), .A2(\mem[16][1] ), .B1(n769), .B2(\mem[18][1] ), 
        .ZN(n513) );
  AOI22D0 U1421 ( .A1(n772), .A2(\mem[17][1] ), .B1(n771), .B2(\mem[19][1] ), 
        .ZN(n512) );
  AOI22D0 U1422 ( .A1(n776), .A2(\mem[25][1] ), .B1(n775), .B2(\mem[27][1] ), 
        .ZN(n510) );
  ND4D0 U1423 ( .A1(n513), .A2(n512), .A3(n511), .A4(n510), .ZN(n519) );
  AOI22D0 U1424 ( .A1(n782), .A2(\mem[20][1] ), .B1(n781), .B2(\mem[22][1] ), 
        .ZN(n517) );
  AOI22D0 U1425 ( .A1(n784), .A2(\mem[21][1] ), .B1(n783), .B2(\mem[23][1] ), 
        .ZN(n516) );
  AOI22D0 U1426 ( .A1(n786), .A2(\mem[28][1] ), .B1(n785), .B2(\mem[29][1] ), 
        .ZN(n515) );
  AOI22D0 U1427 ( .A1(n788), .A2(\mem[31][1] ), .B1(n787), .B2(\mem[0][1] ), 
        .ZN(n514) );
  ND4D0 U1428 ( .A1(n517), .A2(n516), .A3(n515), .A4(n514), .ZN(n518) );
  NR3D0 U1429 ( .A1(n520), .A2(n519), .A3(n518), .ZN(n521) );
  ND4D0 U1430 ( .A1(n524), .A2(n523), .A3(n522), .A4(n521), .ZN(B[1]) );
  AOI22D0 U1431 ( .A1(n746), .A2(\mem[30][4] ), .B1(n745), .B2(\mem[2][4] ), 
        .ZN(n546) );
  AOI22D0 U1432 ( .A1(n748), .A2(\mem[1][4] ), .B1(n747), .B2(\mem[3][4] ), 
        .ZN(n545) );
  AOI22D0 U1433 ( .A1(n750), .A2(\mem[8][4] ), .B1(n749), .B2(\mem[10][4] ), 
        .ZN(n526) );
  AOI22D0 U1434 ( .A1(n752), .A2(\mem[6][4] ), .B1(n751), .B2(\mem[9][4] ), 
        .ZN(n525) );
  OA211D0 U1435 ( .A1(n756), .A2(n527), .B(n526), .C(n525), .Z(n544) );
  AOI22D0 U1436 ( .A1(n758), .A2(\mem[11][4] ), .B1(n757), .B2(\mem[4][4] ), 
        .ZN(n531) );
  AOI22D0 U1437 ( .A1(n760), .A2(\mem[5][4] ), .B1(n759), .B2(\mem[7][4] ), 
        .ZN(n530) );
  AOI22D0 U1438 ( .A1(n762), .A2(\mem[12][4] ), .B1(n761), .B2(\mem[14][4] ), 
        .ZN(n529) );
  AOI22D0 U1439 ( .A1(n764), .A2(\mem[13][4] ), .B1(n763), .B2(\mem[15][4] ), 
        .ZN(n528) );
  ND4D0 U1440 ( .A1(n531), .A2(n530), .A3(n529), .A4(n528), .ZN(n542) );
  AOI22D0 U1441 ( .A1(n770), .A2(\mem[16][4] ), .B1(n769), .B2(\mem[18][4] ), 
        .ZN(n535) );
  AOI22D0 U1442 ( .A1(n772), .A2(\mem[17][4] ), .B1(n771), .B2(\mem[19][4] ), 
        .ZN(n534) );
  AOI22D0 U1443 ( .A1(n774), .A2(\mem[24][4] ), .B1(n773), .B2(\mem[26][4] ), 
        .ZN(n533) );
  AOI22D0 U1444 ( .A1(n776), .A2(\mem[25][4] ), .B1(n775), .B2(\mem[27][4] ), 
        .ZN(n532) );
  ND4D0 U1445 ( .A1(n535), .A2(n534), .A3(n533), .A4(n532), .ZN(n541) );
  AOI22D0 U1446 ( .A1(n782), .A2(\mem[20][4] ), .B1(n781), .B2(\mem[22][4] ), 
        .ZN(n539) );
  AOI22D0 U1447 ( .A1(n784), .A2(\mem[21][4] ), .B1(n783), .B2(\mem[23][4] ), 
        .ZN(n538) );
  AOI22D0 U1448 ( .A1(n786), .A2(\mem[28][4] ), .B1(n785), .B2(\mem[29][4] ), 
        .ZN(n537) );
  AOI22D0 U1449 ( .A1(n788), .A2(\mem[31][4] ), .B1(n787), .B2(\mem[0][4] ), 
        .ZN(n536) );
  ND4D0 U1450 ( .A1(n539), .A2(n538), .A3(n537), .A4(n536), .ZN(n540) );
  NR3D0 U1451 ( .A1(n542), .A2(n541), .A3(n540), .ZN(n543) );
  ND4D0 U1452 ( .A1(n546), .A2(n545), .A3(n544), .A4(n543), .ZN(B[4]) );
  AOI22D0 U1453 ( .A1(n746), .A2(\mem[30][6] ), .B1(n745), .B2(\mem[2][6] ), 
        .ZN(n568) );
  AOI22D0 U1454 ( .A1(n750), .A2(\mem[8][6] ), .B1(n749), .B2(\mem[10][6] ), 
        .ZN(n548) );
  AOI22D0 U1455 ( .A1(n752), .A2(\mem[6][6] ), .B1(n751), .B2(\mem[9][6] ), 
        .ZN(n547) );
  OA211D0 U1456 ( .A1(n756), .A2(n549), .B(n548), .C(n547), .Z(n566) );
  AOI22D0 U1457 ( .A1(n758), .A2(\mem[11][6] ), .B1(n757), .B2(\mem[4][6] ), 
        .ZN(n553) );
  AOI22D0 U1458 ( .A1(n760), .A2(\mem[5][6] ), .B1(n759), .B2(\mem[7][6] ), 
        .ZN(n552) );
  AOI22D0 U1459 ( .A1(n762), .A2(\mem[12][6] ), .B1(n761), .B2(\mem[14][6] ), 
        .ZN(n551) );
  AOI22D0 U1460 ( .A1(n764), .A2(\mem[13][6] ), .B1(n763), .B2(\mem[15][6] ), 
        .ZN(n550) );
  ND4D0 U1461 ( .A1(n553), .A2(n552), .A3(n551), .A4(n550), .ZN(n564) );
  AOI22D0 U1462 ( .A1(n770), .A2(\mem[16][6] ), .B1(n769), .B2(\mem[18][6] ), 
        .ZN(n557) );
  AOI22D0 U1463 ( .A1(n772), .A2(\mem[17][6] ), .B1(n771), .B2(\mem[19][6] ), 
        .ZN(n556) );
  AOI22D0 U1464 ( .A1(n776), .A2(\mem[25][6] ), .B1(n775), .B2(\mem[27][6] ), 
        .ZN(n554) );
  ND4D0 U1465 ( .A1(n557), .A2(n556), .A3(n555), .A4(n554), .ZN(n563) );
  AOI22D0 U1466 ( .A1(n782), .A2(\mem[20][6] ), .B1(n781), .B2(\mem[22][6] ), 
        .ZN(n561) );
  AOI22D0 U1467 ( .A1(n784), .A2(\mem[21][6] ), .B1(n783), .B2(\mem[23][6] ), 
        .ZN(n560) );
  AOI22D0 U1468 ( .A1(n786), .A2(\mem[28][6] ), .B1(n785), .B2(\mem[29][6] ), 
        .ZN(n559) );
  AOI22D0 U1469 ( .A1(n788), .A2(\mem[31][6] ), .B1(n787), .B2(\mem[0][6] ), 
        .ZN(n558) );
  NR3D0 U1470 ( .A1(n564), .A2(n563), .A3(n562), .ZN(n565) );
  ND4D0 U1471 ( .A1(n568), .A2(n567), .A3(n566), .A4(n565), .ZN(B[6]) );
  AOI22D0 U1472 ( .A1(n746), .A2(\mem[30][8] ), .B1(n745), .B2(\mem[2][8] ), 
        .ZN(n590) );
  AOI22D0 U1473 ( .A1(n748), .A2(\mem[1][8] ), .B1(n747), .B2(\mem[3][8] ), 
        .ZN(n589) );
  AOI22D0 U1474 ( .A1(n750), .A2(\mem[8][8] ), .B1(n749), .B2(\mem[10][8] ), 
        .ZN(n570) );
  AOI22D0 U1475 ( .A1(n752), .A2(\mem[6][8] ), .B1(n751), .B2(\mem[9][8] ), 
        .ZN(n569) );
  OA211D0 U1476 ( .A1(n756), .A2(n571), .B(n570), .C(n569), .Z(n588) );
  AOI22D0 U1477 ( .A1(n760), .A2(\mem[5][8] ), .B1(n759), .B2(\mem[7][8] ), 
        .ZN(n574) );
  AOI22D0 U1478 ( .A1(n762), .A2(\mem[12][8] ), .B1(n761), .B2(\mem[14][8] ), 
        .ZN(n573) );
  AOI22D0 U1479 ( .A1(n764), .A2(\mem[13][8] ), .B1(n763), .B2(\mem[15][8] ), 
        .ZN(n572) );
  ND4D0 U1480 ( .A1(n575), .A2(n574), .A3(n573), .A4(n572), .ZN(n586) );
  AOI22D0 U1481 ( .A1(n770), .A2(\mem[16][8] ), .B1(n769), .B2(\mem[18][8] ), 
        .ZN(n579) );
  AOI22D0 U1482 ( .A1(n772), .A2(\mem[17][8] ), .B1(n771), .B2(\mem[19][8] ), 
        .ZN(n578) );
  AOI22D0 U1483 ( .A1(n774), .A2(\mem[24][8] ), .B1(n773), .B2(\mem[26][8] ), 
        .ZN(n577) );
  AOI22D0 U1484 ( .A1(n776), .A2(\mem[25][8] ), .B1(n775), .B2(\mem[27][8] ), 
        .ZN(n576) );
  ND4D0 U1485 ( .A1(n579), .A2(n578), .A3(n577), .A4(n576), .ZN(n585) );
  AOI22D0 U1486 ( .A1(n782), .A2(\mem[20][8] ), .B1(n781), .B2(\mem[22][8] ), 
        .ZN(n583) );
  AOI22D0 U1487 ( .A1(n784), .A2(\mem[21][8] ), .B1(n783), .B2(\mem[23][8] ), 
        .ZN(n582) );
  AOI22D0 U1488 ( .A1(n786), .A2(\mem[28][8] ), .B1(n785), .B2(\mem[29][8] ), 
        .ZN(n581) );
  AOI22D0 U1489 ( .A1(n788), .A2(\mem[31][8] ), .B1(n787), .B2(\mem[0][8] ), 
        .ZN(n580) );
  ND4D0 U1490 ( .A1(n583), .A2(n582), .A3(n581), .A4(n580), .ZN(n584) );
  NR3D0 U1491 ( .A1(n586), .A2(n585), .A3(n584), .ZN(n587) );
  ND4D0 U1492 ( .A1(n590), .A2(n589), .A3(n588), .A4(n587), .ZN(B[8]) );
  AOI22D0 U1493 ( .A1(n746), .A2(\mem[30][10] ), .B1(n745), .B2(\mem[2][10] ), 
        .ZN(n612) );
  AOI22D0 U1494 ( .A1(n748), .A2(\mem[1][10] ), .B1(n747), .B2(\mem[3][10] ), 
        .ZN(n611) );
  AOI22D0 U1495 ( .A1(n750), .A2(\mem[8][10] ), .B1(n749), .B2(\mem[10][10] ), 
        .ZN(n592) );
  AOI22D0 U1496 ( .A1(n752), .A2(\mem[6][10] ), .B1(n751), .B2(\mem[9][10] ), 
        .ZN(n591) );
  AOI22D0 U1497 ( .A1(n758), .A2(\mem[11][10] ), .B1(n757), .B2(\mem[4][10] ), 
        .ZN(n597) );
  AOI22D0 U1498 ( .A1(n760), .A2(\mem[5][10] ), .B1(n759), .B2(\mem[7][10] ), 
        .ZN(n596) );
  AOI22D0 U1499 ( .A1(n762), .A2(\mem[12][10] ), .B1(n761), .B2(\mem[14][10] ), 
        .ZN(n595) );
  AOI22D0 U1500 ( .A1(n764), .A2(\mem[13][10] ), .B1(n763), .B2(\mem[15][10] ), 
        .ZN(n594) );
  ND4D0 U1501 ( .A1(n597), .A2(n596), .A3(n595), .A4(n594), .ZN(n608) );
  AOI22D0 U1502 ( .A1(n770), .A2(\mem[16][10] ), .B1(n769), .B2(\mem[18][10] ), 
        .ZN(n601) );
  AOI22D0 U1503 ( .A1(n772), .A2(\mem[17][10] ), .B1(n771), .B2(\mem[19][10] ), 
        .ZN(n600) );
  AOI22D0 U1504 ( .A1(n774), .A2(\mem[24][10] ), .B1(n773), .B2(\mem[26][10] ), 
        .ZN(n599) );
  AOI22D0 U1505 ( .A1(n776), .A2(\mem[25][10] ), .B1(n775), .B2(\mem[27][10] ), 
        .ZN(n598) );
  ND4D0 U1506 ( .A1(n601), .A2(n600), .A3(n599), .A4(n598), .ZN(n607) );
  AOI22D0 U1507 ( .A1(n782), .A2(\mem[20][10] ), .B1(n781), .B2(\mem[22][10] ), 
        .ZN(n605) );
  AOI22D0 U1508 ( .A1(n786), .A2(\mem[28][10] ), .B1(n785), .B2(\mem[29][10] ), 
        .ZN(n603) );
  AOI22D0 U1509 ( .A1(n788), .A2(\mem[31][10] ), .B1(n787), .B2(\mem[0][10] ), 
        .ZN(n602) );
  ND4D0 U1510 ( .A1(n605), .A2(n604), .A3(n603), .A4(n602), .ZN(n606) );
  NR3D0 U1511 ( .A1(n608), .A2(n607), .A3(n606), .ZN(n609) );
  ND4D0 U1512 ( .A1(n612), .A2(n611), .A3(n610), .A4(n609), .ZN(B[10]) );
  AOI22D0 U1513 ( .A1(n746), .A2(\mem[30][12] ), .B1(n745), .B2(\mem[2][12] ), 
        .ZN(n634) );
  AOI22D0 U1514 ( .A1(n748), .A2(\mem[1][12] ), .B1(n747), .B2(\mem[3][12] ), 
        .ZN(n633) );
  AOI22D0 U1515 ( .A1(n750), .A2(\mem[8][12] ), .B1(n749), .B2(\mem[10][12] ), 
        .ZN(n614) );
  AOI22D0 U1516 ( .A1(n752), .A2(\mem[6][12] ), .B1(n751), .B2(\mem[9][12] ), 
        .ZN(n613) );
  OA211D0 U1517 ( .A1(n756), .A2(n615), .B(n614), .C(n613), .Z(n632) );
  AOI22D0 U1518 ( .A1(n758), .A2(\mem[11][12] ), .B1(n757), .B2(\mem[4][12] ), 
        .ZN(n619) );
  AOI22D0 U1519 ( .A1(n760), .A2(\mem[5][12] ), .B1(n759), .B2(\mem[7][12] ), 
        .ZN(n618) );
  AOI22D0 U1520 ( .A1(n762), .A2(\mem[12][12] ), .B1(n761), .B2(\mem[14][12] ), 
        .ZN(n617) );
  ND4D0 U1521 ( .A1(n619), .A2(n618), .A3(n617), .A4(n616), .ZN(n630) );
  AOI22D0 U1522 ( .A1(n770), .A2(\mem[16][12] ), .B1(n769), .B2(\mem[18][12] ), 
        .ZN(n623) );
  AOI22D0 U1523 ( .A1(n772), .A2(\mem[17][12] ), .B1(n771), .B2(\mem[19][12] ), 
        .ZN(n622) );
  AOI22D0 U1524 ( .A1(n774), .A2(\mem[24][12] ), .B1(n773), .B2(\mem[26][12] ), 
        .ZN(n621) );
  AOI22D0 U1525 ( .A1(n776), .A2(\mem[25][12] ), .B1(n775), .B2(\mem[27][12] ), 
        .ZN(n620) );
  ND4D0 U1526 ( .A1(n623), .A2(n622), .A3(n621), .A4(n620), .ZN(n629) );
  AOI22D0 U1527 ( .A1(n782), .A2(\mem[20][12] ), .B1(n781), .B2(\mem[22][12] ), 
        .ZN(n627) );
  AOI22D0 U1528 ( .A1(n784), .A2(\mem[21][12] ), .B1(n783), .B2(\mem[23][12] ), 
        .ZN(n626) );
  AOI22D0 U1529 ( .A1(n786), .A2(\mem[28][12] ), .B1(n785), .B2(\mem[29][12] ), 
        .ZN(n625) );
  AOI22D0 U1530 ( .A1(n788), .A2(\mem[31][12] ), .B1(n787), .B2(\mem[0][12] ), 
        .ZN(n624) );
  NR3D0 U1531 ( .A1(n630), .A2(n629), .A3(n628), .ZN(n631) );
  ND4D0 U1532 ( .A1(n634), .A2(n633), .A3(n632), .A4(n631), .ZN(B[12]) );
  AOI22D0 U1533 ( .A1(n746), .A2(\mem[30][14] ), .B1(n745), .B2(\mem[2][14] ), 
        .ZN(n656) );
  AOI22D0 U1534 ( .A1(n748), .A2(\mem[1][14] ), .B1(n747), .B2(\mem[3][14] ), 
        .ZN(n655) );
  AOI22D0 U1535 ( .A1(n750), .A2(\mem[8][14] ), .B1(n749), .B2(\mem[10][14] ), 
        .ZN(n636) );
  AOI22D0 U1536 ( .A1(n752), .A2(\mem[6][14] ), .B1(n751), .B2(\mem[9][14] ), 
        .ZN(n635) );
  AOI22D0 U1537 ( .A1(n758), .A2(\mem[11][14] ), .B1(n757), .B2(\mem[4][14] ), 
        .ZN(n641) );
  AOI22D0 U1538 ( .A1(n760), .A2(\mem[5][14] ), .B1(n759), .B2(\mem[7][14] ), 
        .ZN(n640) );
  AOI22D0 U1539 ( .A1(n762), .A2(\mem[12][14] ), .B1(n761), .B2(\mem[14][14] ), 
        .ZN(n639) );
  AOI22D0 U1540 ( .A1(n764), .A2(\mem[13][14] ), .B1(n763), .B2(\mem[15][14] ), 
        .ZN(n638) );
  ND4D0 U1541 ( .A1(n641), .A2(n640), .A3(n639), .A4(n638), .ZN(n652) );
  AOI22D0 U1542 ( .A1(n770), .A2(\mem[16][14] ), .B1(n769), .B2(\mem[18][14] ), 
        .ZN(n645) );
  AOI22D0 U1543 ( .A1(n772), .A2(\mem[17][14] ), .B1(n771), .B2(\mem[19][14] ), 
        .ZN(n644) );
  AOI22D0 U1544 ( .A1(n774), .A2(\mem[24][14] ), .B1(n773), .B2(\mem[26][14] ), 
        .ZN(n643) );
  AOI22D0 U1545 ( .A1(n776), .A2(\mem[25][14] ), .B1(n775), .B2(\mem[27][14] ), 
        .ZN(n642) );
  ND4D0 U1546 ( .A1(n645), .A2(n644), .A3(n643), .A4(n642), .ZN(n651) );
  AOI22D0 U1547 ( .A1(n782), .A2(\mem[20][14] ), .B1(n781), .B2(\mem[22][14] ), 
        .ZN(n649) );
  AOI22D0 U1548 ( .A1(n784), .A2(\mem[21][14] ), .B1(n783), .B2(\mem[23][14] ), 
        .ZN(n648) );
  AOI22D0 U1549 ( .A1(n786), .A2(\mem[28][14] ), .B1(n785), .B2(\mem[29][14] ), 
        .ZN(n647) );
  AOI22D0 U1550 ( .A1(n788), .A2(\mem[31][14] ), .B1(n787), .B2(\mem[0][14] ), 
        .ZN(n646) );
  ND4D0 U1551 ( .A1(n649), .A2(n648), .A3(n647), .A4(n646), .ZN(n650) );
  NR3D0 U1552 ( .A1(n652), .A2(n651), .A3(n650), .ZN(n653) );
  ND4D0 U1553 ( .A1(n656), .A2(n655), .A3(n654), .A4(n653), .ZN(B[14]) );
  AOI22D0 U1554 ( .A1(n746), .A2(\mem[30][16] ), .B1(n745), .B2(\mem[2][16] ), 
        .ZN(n678) );
  AOI22D0 U1555 ( .A1(n748), .A2(\mem[1][16] ), .B1(n747), .B2(\mem[3][16] ), 
        .ZN(n677) );
  AOI22D0 U1556 ( .A1(n750), .A2(\mem[8][16] ), .B1(n749), .B2(\mem[10][16] ), 
        .ZN(n658) );
  AOI22D0 U1557 ( .A1(n752), .A2(\mem[6][16] ), .B1(n751), .B2(\mem[9][16] ), 
        .ZN(n657) );
  OA211D0 U1558 ( .A1(n756), .A2(n659), .B(n658), .C(n657), .Z(n676) );
  AOI22D0 U1559 ( .A1(n758), .A2(\mem[11][16] ), .B1(n757), .B2(\mem[4][16] ), 
        .ZN(n663) );
  AOI22D0 U1560 ( .A1(n760), .A2(\mem[5][16] ), .B1(n759), .B2(\mem[7][16] ), 
        .ZN(n662) );
  AOI22D0 U1561 ( .A1(n762), .A2(\mem[12][16] ), .B1(n761), .B2(\mem[14][16] ), 
        .ZN(n661) );
  AOI22D0 U1562 ( .A1(n764), .A2(\mem[13][16] ), .B1(n763), .B2(\mem[15][16] ), 
        .ZN(n660) );
  ND4D0 U1563 ( .A1(n663), .A2(n662), .A3(n661), .A4(n660), .ZN(n674) );
  AOI22D0 U1564 ( .A1(n770), .A2(\mem[16][16] ), .B1(n769), .B2(\mem[18][16] ), 
        .ZN(n667) );
  AOI22D0 U1565 ( .A1(n772), .A2(\mem[17][16] ), .B1(n771), .B2(\mem[19][16] ), 
        .ZN(n666) );
  AOI22D0 U1566 ( .A1(n776), .A2(\mem[25][16] ), .B1(n775), .B2(\mem[27][16] ), 
        .ZN(n664) );
  ND4D0 U1567 ( .A1(n667), .A2(n666), .A3(n665), .A4(n664), .ZN(n673) );
  AOI22D0 U1568 ( .A1(n782), .A2(\mem[20][16] ), .B1(n781), .B2(\mem[22][16] ), 
        .ZN(n671) );
  AOI22D0 U1569 ( .A1(n784), .A2(\mem[21][16] ), .B1(n783), .B2(\mem[23][16] ), 
        .ZN(n670) );
  AOI22D0 U1570 ( .A1(n786), .A2(\mem[28][16] ), .B1(n785), .B2(\mem[29][16] ), 
        .ZN(n669) );
  AOI22D0 U1571 ( .A1(n788), .A2(\mem[31][16] ), .B1(n787), .B2(\mem[0][16] ), 
        .ZN(n668) );
  ND4D0 U1572 ( .A1(n671), .A2(n670), .A3(n669), .A4(n668), .ZN(n672) );
  NR3D0 U1573 ( .A1(n674), .A2(n673), .A3(n672), .ZN(n675) );
  ND4D0 U1574 ( .A1(n678), .A2(n677), .A3(n676), .A4(n675), .ZN(B[16]) );
  AOI22D0 U1575 ( .A1(n746), .A2(\mem[30][18] ), .B1(n745), .B2(\mem[2][18] ), 
        .ZN(n700) );
  AOI22D0 U1576 ( .A1(n748), .A2(\mem[1][18] ), .B1(n747), .B2(\mem[3][18] ), 
        .ZN(n699) );
  AOI22D0 U1577 ( .A1(n750), .A2(\mem[8][18] ), .B1(n749), .B2(\mem[10][18] ), 
        .ZN(n680) );
  AOI22D0 U1578 ( .A1(n752), .A2(\mem[6][18] ), .B1(n751), .B2(\mem[9][18] ), 
        .ZN(n679) );
  OA211D0 U1579 ( .A1(n756), .A2(n681), .B(n680), .C(n679), .Z(n698) );
  AOI22D0 U1580 ( .A1(n760), .A2(\mem[5][18] ), .B1(n759), .B2(\mem[7][18] ), 
        .ZN(n684) );
  AOI22D0 U1581 ( .A1(n762), .A2(\mem[12][18] ), .B1(n761), .B2(\mem[14][18] ), 
        .ZN(n683) );
  AOI22D0 U1582 ( .A1(n764), .A2(\mem[13][18] ), .B1(n763), .B2(\mem[15][18] ), 
        .ZN(n682) );
  ND4D0 U1583 ( .A1(n685), .A2(n684), .A3(n683), .A4(n682), .ZN(n696) );
  AOI22D0 U1584 ( .A1(n770), .A2(\mem[16][18] ), .B1(n769), .B2(\mem[18][18] ), 
        .ZN(n689) );
  AOI22D0 U1585 ( .A1(n772), .A2(\mem[17][18] ), .B1(n771), .B2(\mem[19][18] ), 
        .ZN(n688) );
  AOI22D0 U1586 ( .A1(n774), .A2(\mem[24][18] ), .B1(n773), .B2(\mem[26][18] ), 
        .ZN(n687) );
  AOI22D0 U1587 ( .A1(n776), .A2(\mem[25][18] ), .B1(n775), .B2(\mem[27][18] ), 
        .ZN(n686) );
  ND4D0 U1588 ( .A1(n689), .A2(n688), .A3(n687), .A4(n686), .ZN(n695) );
  AOI22D0 U1589 ( .A1(n782), .A2(\mem[20][18] ), .B1(n781), .B2(\mem[22][18] ), 
        .ZN(n693) );
  AOI22D0 U1590 ( .A1(n784), .A2(\mem[21][18] ), .B1(n783), .B2(\mem[23][18] ), 
        .ZN(n692) );
  AOI22D0 U1591 ( .A1(n786), .A2(\mem[28][18] ), .B1(n785), .B2(\mem[29][18] ), 
        .ZN(n691) );
  AOI22D0 U1592 ( .A1(n788), .A2(\mem[31][18] ), .B1(n787), .B2(\mem[0][18] ), 
        .ZN(n690) );
  NR3D0 U1593 ( .A1(n696), .A2(n695), .A3(n694), .ZN(n697) );
  ND4D0 U1594 ( .A1(n700), .A2(n699), .A3(n698), .A4(n697), .ZN(B[18]) );
  AOI22D0 U1595 ( .A1(n746), .A2(\mem[30][20] ), .B1(n745), .B2(\mem[2][20] ), 
        .ZN(n722) );
  AOI22D0 U1596 ( .A1(n748), .A2(\mem[1][20] ), .B1(n747), .B2(\mem[3][20] ), 
        .ZN(n721) );
  AOI22D0 U1597 ( .A1(n750), .A2(\mem[8][20] ), .B1(n749), .B2(\mem[10][20] ), 
        .ZN(n702) );
  AOI22D0 U1598 ( .A1(n752), .A2(\mem[6][20] ), .B1(n751), .B2(\mem[9][20] ), 
        .ZN(n701) );
  OA211D0 U1599 ( .A1(n756), .A2(n703), .B(n702), .C(n701), .Z(n720) );
  AOI22D0 U1600 ( .A1(n758), .A2(\mem[11][20] ), .B1(n757), .B2(\mem[4][20] ), 
        .ZN(n707) );
  AOI22D0 U1601 ( .A1(n760), .A2(\mem[5][20] ), .B1(n759), .B2(\mem[7][20] ), 
        .ZN(n706) );
  AOI22D0 U1602 ( .A1(n762), .A2(\mem[12][20] ), .B1(n761), .B2(\mem[14][20] ), 
        .ZN(n705) );
  AOI22D0 U1603 ( .A1(n764), .A2(\mem[13][20] ), .B1(n763), .B2(\mem[15][20] ), 
        .ZN(n704) );
  ND4D0 U1604 ( .A1(n707), .A2(n706), .A3(n705), .A4(n704), .ZN(n718) );
  AOI22D0 U1605 ( .A1(n770), .A2(\mem[16][20] ), .B1(n769), .B2(\mem[18][20] ), 
        .ZN(n711) );
  AOI22D0 U1606 ( .A1(n772), .A2(\mem[17][20] ), .B1(n771), .B2(\mem[19][20] ), 
        .ZN(n710) );
  AOI22D0 U1607 ( .A1(n774), .A2(\mem[24][20] ), .B1(n773), .B2(\mem[26][20] ), 
        .ZN(n709) );
  AOI22D0 U1608 ( .A1(n776), .A2(\mem[25][20] ), .B1(n775), .B2(\mem[27][20] ), 
        .ZN(n708) );
  ND4D0 U1609 ( .A1(n711), .A2(n710), .A3(n709), .A4(n708), .ZN(n717) );
  AOI22D0 U1610 ( .A1(n782), .A2(\mem[20][20] ), .B1(n781), .B2(\mem[22][20] ), 
        .ZN(n715) );
  AOI22D0 U1611 ( .A1(n786), .A2(\mem[28][20] ), .B1(n785), .B2(\mem[29][20] ), 
        .ZN(n713) );
  AOI22D0 U1612 ( .A1(n788), .A2(\mem[31][20] ), .B1(n787), .B2(\mem[0][20] ), 
        .ZN(n712) );
  ND4D0 U1613 ( .A1(n715), .A2(n714), .A3(n713), .A4(n712), .ZN(n716) );
  NR3D0 U1614 ( .A1(n718), .A2(n717), .A3(n716), .ZN(n719) );
  ND4D0 U1615 ( .A1(n722), .A2(n721), .A3(n720), .A4(n719), .ZN(B[20]) );
  AOI22D0 U1616 ( .A1(n746), .A2(\mem[30][22] ), .B1(n745), .B2(\mem[2][22] ), 
        .ZN(n744) );
  AOI22D0 U1617 ( .A1(n748), .A2(\mem[1][22] ), .B1(n747), .B2(\mem[3][22] ), 
        .ZN(n743) );
  AOI22D0 U1618 ( .A1(n750), .A2(\mem[8][22] ), .B1(n749), .B2(\mem[10][22] ), 
        .ZN(n724) );
  AOI22D0 U1619 ( .A1(n752), .A2(\mem[6][22] ), .B1(n751), .B2(\mem[9][22] ), 
        .ZN(n723) );
  OA211D0 U1620 ( .A1(n756), .A2(n725), .B(n724), .C(n723), .Z(n742) );
  AOI22D0 U1621 ( .A1(n758), .A2(\mem[11][22] ), .B1(n757), .B2(\mem[4][22] ), 
        .ZN(n729) );
  AOI22D0 U1622 ( .A1(n760), .A2(\mem[5][22] ), .B1(n759), .B2(\mem[7][22] ), 
        .ZN(n728) );
  AOI22D0 U1623 ( .A1(n762), .A2(\mem[12][22] ), .B1(n761), .B2(\mem[14][22] ), 
        .ZN(n727) );
  ND4D0 U1624 ( .A1(n729), .A2(n728), .A3(n727), .A4(n726), .ZN(n740) );
  AOI22D0 U1625 ( .A1(n770), .A2(\mem[16][22] ), .B1(n769), .B2(\mem[18][22] ), 
        .ZN(n733) );
  AOI22D0 U1626 ( .A1(n772), .A2(\mem[17][22] ), .B1(n771), .B2(\mem[19][22] ), 
        .ZN(n732) );
  AOI22D0 U1627 ( .A1(n774), .A2(\mem[24][22] ), .B1(n773), .B2(\mem[26][22] ), 
        .ZN(n731) );
  AOI22D0 U1628 ( .A1(n776), .A2(\mem[25][22] ), .B1(n775), .B2(\mem[27][22] ), 
        .ZN(n730) );
  ND4D0 U1629 ( .A1(n733), .A2(n732), .A3(n731), .A4(n730), .ZN(n739) );
  AOI22D0 U1630 ( .A1(n782), .A2(\mem[20][22] ), .B1(n781), .B2(\mem[22][22] ), 
        .ZN(n737) );
  AOI22D0 U1631 ( .A1(n784), .A2(\mem[21][22] ), .B1(n783), .B2(\mem[23][22] ), 
        .ZN(n736) );
  AOI22D0 U1632 ( .A1(n786), .A2(\mem[28][22] ), .B1(n785), .B2(\mem[29][22] ), 
        .ZN(n735) );
  AOI22D0 U1633 ( .A1(n788), .A2(\mem[31][22] ), .B1(n787), .B2(\mem[0][22] ), 
        .ZN(n734) );
  ND4D0 U1634 ( .A1(n737), .A2(n736), .A3(n735), .A4(n734), .ZN(n738) );
  NR3D0 U1635 ( .A1(n740), .A2(n739), .A3(n738), .ZN(n741) );
  AOI22D0 U1636 ( .A1(n748), .A2(\mem[1][2] ), .B1(n747), .B2(\mem[3][2] ), 
        .ZN(n798) );
  AOI22D0 U1637 ( .A1(n750), .A2(\mem[8][2] ), .B1(n749), .B2(\mem[10][2] ), 
        .ZN(n754) );
  AOI22D0 U1638 ( .A1(n752), .A2(\mem[6][2] ), .B1(n751), .B2(\mem[9][2] ), 
        .ZN(n753) );
  OA211D0 U1639 ( .A1(n756), .A2(n755), .B(n754), .C(n753), .Z(n797) );
  AOI22D0 U1640 ( .A1(n758), .A2(\mem[11][2] ), .B1(n757), .B2(\mem[4][2] ), 
        .ZN(n768) );
  AOI22D0 U1641 ( .A1(n760), .A2(\mem[5][2] ), .B1(n759), .B2(\mem[7][2] ), 
        .ZN(n767) );
  AOI22D0 U1642 ( .A1(n762), .A2(\mem[12][2] ), .B1(n761), .B2(\mem[14][2] ), 
        .ZN(n766) );
  ND4D0 U1643 ( .A1(n768), .A2(n767), .A3(n766), .A4(n765), .ZN(n795) );
  AOI22D0 U1644 ( .A1(n770), .A2(\mem[16][2] ), .B1(n769), .B2(\mem[18][2] ), 
        .ZN(n780) );
  AOI22D0 U1645 ( .A1(n772), .A2(\mem[17][2] ), .B1(n771), .B2(\mem[19][2] ), 
        .ZN(n779) );
  AOI22D0 U1646 ( .A1(n774), .A2(\mem[24][2] ), .B1(n773), .B2(\mem[26][2] ), 
        .ZN(n778) );
  AOI22D0 U1647 ( .A1(n776), .A2(\mem[25][2] ), .B1(n775), .B2(\mem[27][2] ), 
        .ZN(n777) );
  ND4D0 U1648 ( .A1(n780), .A2(n779), .A3(n778), .A4(n777), .ZN(n794) );
  AOI22D0 U1649 ( .A1(n782), .A2(\mem[20][2] ), .B1(n781), .B2(\mem[22][2] ), 
        .ZN(n792) );
  AOI22D0 U1650 ( .A1(n784), .A2(\mem[21][2] ), .B1(n783), .B2(\mem[23][2] ), 
        .ZN(n791) );
  AOI22D0 U1651 ( .A1(n786), .A2(\mem[28][2] ), .B1(n785), .B2(\mem[29][2] ), 
        .ZN(n790) );
  AOI22D0 U1652 ( .A1(n788), .A2(\mem[31][2] ), .B1(n787), .B2(\mem[0][2] ), 
        .ZN(n789) );
  ND4D0 U1653 ( .A1(n792), .A2(n791), .A3(n790), .A4(n789), .ZN(n793) );
  NR3D0 U1654 ( .A1(n795), .A2(n794), .A3(n793), .ZN(n796) );
  ND4D0 U1655 ( .A1(n799), .A2(n798), .A3(n797), .A4(n796), .ZN(B[2]) );
  AOI22D0 U1656 ( .A1(\mem[0][23] ), .A2(n1121), .B1(\mem[2][23] ), .B2(n1120), 
        .ZN(n803) );
  AOI22D0 U1657 ( .A1(\mem[1][23] ), .A2(n1123), .B1(\mem[3][23] ), .B2(n1122), 
        .ZN(n802) );
  AOI22D0 U1658 ( .A1(\mem[8][23] ), .A2(n1125), .B1(\mem[10][23] ), .B2(n1124), .ZN(n801) );
  AOI22D0 U1659 ( .A1(\mem[11][23] ), .A2(n1127), .B1(\mem[9][23] ), .B2(n1126), .ZN(n800) );
  ND4D0 U1660 ( .A1(n803), .A2(n802), .A3(n801), .A4(n800), .ZN(n819) );
  AOI22D0 U1661 ( .A1(\mem[4][23] ), .A2(n1133), .B1(\mem[6][23] ), .B2(n1132), 
        .ZN(n807) );
  AOI22D0 U1662 ( .A1(\mem[5][23] ), .A2(n1135), .B1(\mem[7][23] ), .B2(n1134), 
        .ZN(n806) );
  AOI22D0 U1663 ( .A1(\mem[12][23] ), .A2(n1137), .B1(\mem[14][23] ), .B2(
        n1136), .ZN(n805) );
  AOI22D0 U1664 ( .A1(\mem[13][23] ), .A2(n1139), .B1(\mem[15][23] ), .B2(
        n1138), .ZN(n804) );
  AOI22D0 U1665 ( .A1(\mem[17][23] ), .A2(n1147), .B1(\mem[19][23] ), .B2(
        n1146), .ZN(n810) );
  AOI22D0 U1666 ( .A1(\mem[24][23] ), .A2(n1149), .B1(\mem[26][23] ), .B2(
        n1148), .ZN(n809) );
  AOI22D0 U1667 ( .A1(\mem[25][23] ), .A2(n1151), .B1(\mem[27][23] ), .B2(
        n1150), .ZN(n808) );
  ND4D0 U1668 ( .A1(n811), .A2(n810), .A3(n809), .A4(n808), .ZN(n817) );
  AOI22D0 U1669 ( .A1(\mem[20][23] ), .A2(n1157), .B1(\mem[22][23] ), .B2(
        n1156), .ZN(n815) );
  AOI22D0 U1670 ( .A1(\mem[21][23] ), .A2(n1159), .B1(\mem[23][23] ), .B2(
        n1158), .ZN(n814) );
  AOI22D0 U1671 ( .A1(\mem[28][23] ), .A2(n1161), .B1(\mem[30][23] ), .B2(
        n1160), .ZN(n813) );
  AOI22D0 U1672 ( .A1(\mem[29][23] ), .A2(n1163), .B1(\mem[31][23] ), .B2(
        n1162), .ZN(n812) );
  ND4D0 U1673 ( .A1(n815), .A2(n814), .A3(n813), .A4(n812), .ZN(n816) );
  OR4D0 U1674 ( .A1(n819), .A2(n818), .A3(n817), .A4(n816), .Z(A[23]) );
  AOI22D0 U1675 ( .A1(\mem[0][22] ), .A2(n1121), .B1(\mem[2][22] ), .B2(n1120), 
        .ZN(n823) );
  AOI22D0 U1676 ( .A1(\mem[1][22] ), .A2(n1123), .B1(\mem[3][22] ), .B2(n1122), 
        .ZN(n822) );
  AOI22D0 U1677 ( .A1(\mem[8][22] ), .A2(n1125), .B1(\mem[10][22] ), .B2(n1124), .ZN(n821) );
  AOI22D0 U1678 ( .A1(\mem[11][22] ), .A2(n1127), .B1(\mem[9][22] ), .B2(n1126), .ZN(n820) );
  ND4D0 U1679 ( .A1(n823), .A2(n822), .A3(n821), .A4(n820), .ZN(n839) );
  AOI22D0 U1680 ( .A1(\mem[4][22] ), .A2(n1133), .B1(\mem[6][22] ), .B2(n1132), 
        .ZN(n827) );
  AOI22D0 U1681 ( .A1(\mem[5][22] ), .A2(n1135), .B1(\mem[7][22] ), .B2(n1134), 
        .ZN(n826) );
  AOI22D0 U1682 ( .A1(\mem[12][22] ), .A2(n1137), .B1(\mem[14][22] ), .B2(
        n1136), .ZN(n825) );
  ND4D0 U1683 ( .A1(n827), .A2(n826), .A3(n825), .A4(n824), .ZN(n838) );
  AOI22D0 U1684 ( .A1(\mem[16][22] ), .A2(n1145), .B1(\mem[18][22] ), .B2(
        n1144), .ZN(n831) );
  AOI22D0 U1685 ( .A1(\mem[17][22] ), .A2(n1147), .B1(\mem[19][22] ), .B2(
        n1146), .ZN(n830) );
  AOI22D0 U1686 ( .A1(\mem[24][22] ), .A2(n1149), .B1(\mem[26][22] ), .B2(
        n1148), .ZN(n829) );
  AOI22D0 U1687 ( .A1(\mem[25][22] ), .A2(n1151), .B1(\mem[27][22] ), .B2(
        n1150), .ZN(n828) );
  ND4D0 U1688 ( .A1(n831), .A2(n830), .A3(n829), .A4(n828), .ZN(n837) );
  AOI22D0 U1689 ( .A1(\mem[20][22] ), .A2(n1157), .B1(\mem[22][22] ), .B2(
        n1156), .ZN(n835) );
  AOI22D0 U1690 ( .A1(\mem[21][22] ), .A2(n1159), .B1(\mem[23][22] ), .B2(
        n1158), .ZN(n834) );
  AOI22D0 U1691 ( .A1(\mem[28][22] ), .A2(n1161), .B1(\mem[30][22] ), .B2(
        n1160), .ZN(n833) );
  AOI22D0 U1692 ( .A1(\mem[29][22] ), .A2(n1163), .B1(\mem[31][22] ), .B2(
        n1162), .ZN(n832) );
  ND4D0 U1693 ( .A1(n835), .A2(n834), .A3(n833), .A4(n832), .ZN(n836) );
  OR4D0 U1694 ( .A1(n839), .A2(n838), .A3(n837), .A4(n836), .Z(A[22]) );
  AOI22D0 U1695 ( .A1(\mem[0][19] ), .A2(n1121), .B1(\mem[2][19] ), .B2(n1120), 
        .ZN(n843) );
  AOI22D0 U1696 ( .A1(\mem[1][19] ), .A2(n1123), .B1(\mem[3][19] ), .B2(n1122), 
        .ZN(n842) );
  AOI22D0 U1697 ( .A1(\mem[8][19] ), .A2(n1125), .B1(\mem[10][19] ), .B2(n1124), .ZN(n841) );
  AOI22D0 U1698 ( .A1(\mem[11][19] ), .A2(n1127), .B1(\mem[9][19] ), .B2(n1126), .ZN(n840) );
  AOI22D0 U1699 ( .A1(\mem[5][19] ), .A2(n1135), .B1(\mem[7][19] ), .B2(n1134), 
        .ZN(n846) );
  AOI22D0 U1700 ( .A1(\mem[12][19] ), .A2(n1137), .B1(\mem[14][19] ), .B2(
        n1136), .ZN(n845) );
  AOI22D0 U1701 ( .A1(\mem[13][19] ), .A2(n1139), .B1(\mem[15][19] ), .B2(
        n1138), .ZN(n844) );
  ND4D0 U1702 ( .A1(n847), .A2(n846), .A3(n845), .A4(n844), .ZN(n858) );
  AOI22D0 U1703 ( .A1(\mem[16][19] ), .A2(n1145), .B1(\mem[18][19] ), .B2(
        n1144), .ZN(n851) );
  AOI22D0 U1704 ( .A1(\mem[17][19] ), .A2(n1147), .B1(\mem[19][19] ), .B2(
        n1146), .ZN(n850) );
  AOI22D0 U1705 ( .A1(\mem[24][19] ), .A2(n1149), .B1(\mem[26][19] ), .B2(
        n1148), .ZN(n849) );
  AOI22D0 U1706 ( .A1(\mem[25][19] ), .A2(n1151), .B1(\mem[27][19] ), .B2(
        n1150), .ZN(n848) );
  ND4D0 U1707 ( .A1(n851), .A2(n850), .A3(n849), .A4(n848), .ZN(n857) );
  AOI22D0 U1708 ( .A1(\mem[20][19] ), .A2(n1157), .B1(\mem[22][19] ), .B2(
        n1156), .ZN(n855) );
  AOI22D0 U1709 ( .A1(\mem[21][19] ), .A2(n1159), .B1(\mem[23][19] ), .B2(
        n1158), .ZN(n854) );
  AOI22D0 U1710 ( .A1(\mem[28][19] ), .A2(n1161), .B1(\mem[30][19] ), .B2(
        n1160), .ZN(n853) );
  AOI22D0 U1711 ( .A1(\mem[29][19] ), .A2(n1163), .B1(\mem[31][19] ), .B2(
        n1162), .ZN(n852) );
  ND4D0 U1712 ( .A1(n855), .A2(n854), .A3(n853), .A4(n852), .ZN(n856) );
  OR4D0 U1713 ( .A1(n859), .A2(n858), .A3(n857), .A4(n856), .Z(A[19]) );
  AOI22D0 U1714 ( .A1(\mem[0][18] ), .A2(n1121), .B1(\mem[2][18] ), .B2(n1120), 
        .ZN(n863) );
  AOI22D0 U1715 ( .A1(\mem[1][18] ), .A2(n1123), .B1(\mem[3][18] ), .B2(n1122), 
        .ZN(n862) );
  AOI22D0 U1716 ( .A1(\mem[8][18] ), .A2(n1125), .B1(\mem[10][18] ), .B2(n1124), .ZN(n861) );
  ND4D0 U1717 ( .A1(n863), .A2(n862), .A3(n861), .A4(n860), .ZN(n879) );
  AOI22D0 U1718 ( .A1(\mem[4][18] ), .A2(n1133), .B1(\mem[6][18] ), .B2(n1132), 
        .ZN(n867) );
  AOI22D0 U1719 ( .A1(\mem[5][18] ), .A2(n1135), .B1(\mem[7][18] ), .B2(n1134), 
        .ZN(n866) );
  AOI22D0 U1720 ( .A1(\mem[12][18] ), .A2(n1137), .B1(\mem[14][18] ), .B2(
        n1136), .ZN(n865) );
  AOI22D0 U1721 ( .A1(\mem[13][18] ), .A2(n1139), .B1(\mem[15][18] ), .B2(
        n1138), .ZN(n864) );
  ND4D0 U1722 ( .A1(n867), .A2(n866), .A3(n865), .A4(n864), .ZN(n878) );
  AOI22D0 U1723 ( .A1(\mem[16][18] ), .A2(n1145), .B1(\mem[18][18] ), .B2(
        n1144), .ZN(n871) );
  AOI22D0 U1724 ( .A1(\mem[17][18] ), .A2(n1147), .B1(\mem[19][18] ), .B2(
        n1146), .ZN(n870) );
  AOI22D0 U1725 ( .A1(\mem[24][18] ), .A2(n1149), .B1(\mem[26][18] ), .B2(
        n1148), .ZN(n869) );
  AOI22D0 U1726 ( .A1(\mem[25][18] ), .A2(n1151), .B1(\mem[27][18] ), .B2(
        n1150), .ZN(n868) );
  ND4D0 U1727 ( .A1(n871), .A2(n870), .A3(n869), .A4(n868), .ZN(n877) );
  AOI22D0 U1728 ( .A1(\mem[20][18] ), .A2(n1157), .B1(\mem[22][18] ), .B2(
        n1156), .ZN(n875) );
  AOI22D0 U1729 ( .A1(\mem[21][18] ), .A2(n1159), .B1(\mem[23][18] ), .B2(
        n1158), .ZN(n874) );
  AOI22D0 U1730 ( .A1(\mem[28][18] ), .A2(n1161), .B1(\mem[30][18] ), .B2(
        n1160), .ZN(n873) );
  AOI22D0 U1731 ( .A1(\mem[29][18] ), .A2(n1163), .B1(\mem[31][18] ), .B2(
        n1162), .ZN(n872) );
  ND4D0 U1732 ( .A1(n875), .A2(n874), .A3(n873), .A4(n872), .ZN(n876) );
  OR4D0 U1733 ( .A1(n879), .A2(n878), .A3(n877), .A4(n876), .Z(A[18]) );
  AOI22D0 U1734 ( .A1(\mem[0][16] ), .A2(n1121), .B1(\mem[2][16] ), .B2(n1120), 
        .ZN(n883) );
  AOI22D0 U1735 ( .A1(\mem[8][16] ), .A2(n1125), .B1(\mem[10][16] ), .B2(n1124), .ZN(n881) );
  AOI22D0 U1736 ( .A1(\mem[11][16] ), .A2(n1127), .B1(\mem[9][16] ), .B2(n1126), .ZN(n880) );
  ND4D0 U1737 ( .A1(n883), .A2(n882), .A3(n881), .A4(n880), .ZN(n899) );
  AOI22D0 U1738 ( .A1(\mem[4][16] ), .A2(n1133), .B1(\mem[6][16] ), .B2(n1132), 
        .ZN(n887) );
  AOI22D0 U1739 ( .A1(\mem[5][16] ), .A2(n1135), .B1(\mem[7][16] ), .B2(n1134), 
        .ZN(n886) );
  AOI22D0 U1740 ( .A1(\mem[12][16] ), .A2(n1137), .B1(\mem[14][16] ), .B2(
        n1136), .ZN(n885) );
  AOI22D0 U1741 ( .A1(\mem[13][16] ), .A2(n1139), .B1(\mem[15][16] ), .B2(
        n1138), .ZN(n884) );
  ND4D0 U1742 ( .A1(n887), .A2(n886), .A3(n885), .A4(n884), .ZN(n898) );
  AOI22D0 U1743 ( .A1(\mem[16][16] ), .A2(n1145), .B1(\mem[18][16] ), .B2(
        n1144), .ZN(n891) );
  AOI22D0 U1744 ( .A1(\mem[17][16] ), .A2(n1147), .B1(\mem[19][16] ), .B2(
        n1146), .ZN(n890) );
  AOI22D0 U1745 ( .A1(\mem[24][16] ), .A2(n1149), .B1(\mem[26][16] ), .B2(
        n1148), .ZN(n889) );
  AOI22D0 U1746 ( .A1(\mem[25][16] ), .A2(n1151), .B1(\mem[27][16] ), .B2(
        n1150), .ZN(n888) );
  ND4D0 U1747 ( .A1(n891), .A2(n890), .A3(n889), .A4(n888), .ZN(n897) );
  AOI22D0 U1748 ( .A1(\mem[20][16] ), .A2(n1157), .B1(\mem[22][16] ), .B2(
        n1156), .ZN(n895) );
  AOI22D0 U1749 ( .A1(\mem[21][16] ), .A2(n1159), .B1(\mem[23][16] ), .B2(
        n1158), .ZN(n894) );
  AOI22D0 U1750 ( .A1(\mem[28][16] ), .A2(n1161), .B1(\mem[30][16] ), .B2(
        n1160), .ZN(n893) );
  AOI22D0 U1751 ( .A1(\mem[29][16] ), .A2(n1163), .B1(\mem[31][16] ), .B2(
        n1162), .ZN(n892) );
  OR4D0 U1752 ( .A1(n899), .A2(n898), .A3(n897), .A4(n896), .Z(A[16]) );
  AOI22D0 U1753 ( .A1(\mem[0][13] ), .A2(n1121), .B1(\mem[2][13] ), .B2(n1120), 
        .ZN(n903) );
  AOI22D0 U1754 ( .A1(\mem[1][13] ), .A2(n1123), .B1(\mem[3][13] ), .B2(n1122), 
        .ZN(n902) );
  AOI22D0 U1755 ( .A1(\mem[8][13] ), .A2(n1125), .B1(\mem[10][13] ), .B2(n1124), .ZN(n901) );
  AOI22D0 U1756 ( .A1(\mem[11][13] ), .A2(n1127), .B1(\mem[9][13] ), .B2(n1126), .ZN(n900) );
  ND4D0 U1757 ( .A1(n903), .A2(n902), .A3(n901), .A4(n900), .ZN(n919) );
  AOI22D0 U1758 ( .A1(\mem[4][13] ), .A2(n1133), .B1(\mem[6][13] ), .B2(n1132), 
        .ZN(n907) );
  AOI22D0 U1759 ( .A1(\mem[5][13] ), .A2(n1135), .B1(\mem[7][13] ), .B2(n1134), 
        .ZN(n906) );
  AOI22D0 U1760 ( .A1(\mem[12][13] ), .A2(n1137), .B1(\mem[14][13] ), .B2(
        n1136), .ZN(n905) );
  AOI22D0 U1761 ( .A1(\mem[13][13] ), .A2(n1139), .B1(\mem[15][13] ), .B2(
        n1138), .ZN(n904) );
  ND4D0 U1762 ( .A1(n907), .A2(n906), .A3(n905), .A4(n904), .ZN(n918) );
  AOI22D0 U1763 ( .A1(\mem[16][13] ), .A2(n1145), .B1(\mem[18][13] ), .B2(
        n1144), .ZN(n911) );
  AOI22D0 U1764 ( .A1(\mem[17][13] ), .A2(n1147), .B1(\mem[19][13] ), .B2(
        n1146), .ZN(n910) );
  AOI22D0 U1765 ( .A1(\mem[24][13] ), .A2(n1149), .B1(\mem[26][13] ), .B2(
        n1148), .ZN(n909) );
  AOI22D0 U1766 ( .A1(\mem[25][13] ), .A2(n1151), .B1(\mem[27][13] ), .B2(
        n1150), .ZN(n908) );
  ND4D0 U1767 ( .A1(n911), .A2(n910), .A3(n909), .A4(n908), .ZN(n917) );
  AOI22D0 U1768 ( .A1(\mem[20][13] ), .A2(n1157), .B1(\mem[22][13] ), .B2(
        n1156), .ZN(n915) );
  AOI22D0 U1769 ( .A1(\mem[28][13] ), .A2(n1161), .B1(\mem[30][13] ), .B2(
        n1160), .ZN(n913) );
  AOI22D0 U1770 ( .A1(\mem[29][13] ), .A2(n1163), .B1(\mem[31][13] ), .B2(
        n1162), .ZN(n912) );
  ND4D0 U1771 ( .A1(n915), .A2(n914), .A3(n913), .A4(n912), .ZN(n916) );
  OR4D0 U1772 ( .A1(n919), .A2(n918), .A3(n917), .A4(n916), .Z(A[13]) );
  AOI22D0 U1773 ( .A1(\mem[0][12] ), .A2(n1121), .B1(\mem[2][12] ), .B2(n1120), 
        .ZN(n923) );
  AOI22D0 U1774 ( .A1(\mem[1][12] ), .A2(n1123), .B1(\mem[3][12] ), .B2(n1122), 
        .ZN(n922) );
  AOI22D0 U1775 ( .A1(\mem[8][12] ), .A2(n1125), .B1(\mem[10][12] ), .B2(n1124), .ZN(n921) );
  AOI22D0 U1776 ( .A1(\mem[11][12] ), .A2(n1127), .B1(\mem[9][12] ), .B2(n1126), .ZN(n920) );
  ND4D0 U1777 ( .A1(n923), .A2(n922), .A3(n921), .A4(n920), .ZN(n939) );
  AOI22D0 U1778 ( .A1(\mem[4][12] ), .A2(n1133), .B1(\mem[6][12] ), .B2(n1132), 
        .ZN(n927) );
  AOI22D0 U1779 ( .A1(\mem[5][12] ), .A2(n1135), .B1(\mem[7][12] ), .B2(n1134), 
        .ZN(n926) );
  AOI22D0 U1780 ( .A1(\mem[12][12] ), .A2(n1137), .B1(\mem[14][12] ), .B2(
        n1136), .ZN(n925) );
  AOI22D0 U1781 ( .A1(\mem[13][12] ), .A2(n1139), .B1(\mem[15][12] ), .B2(
        n1138), .ZN(n924) );
  ND4D0 U1782 ( .A1(n927), .A2(n926), .A3(n925), .A4(n924), .ZN(n938) );
  AOI22D0 U1783 ( .A1(\mem[16][12] ), .A2(n1145), .B1(\mem[18][12] ), .B2(
        n1144), .ZN(n931) );
  AOI22D0 U1784 ( .A1(\mem[17][12] ), .A2(n1147), .B1(\mem[19][12] ), .B2(
        n1146), .ZN(n930) );
  AOI22D0 U1785 ( .A1(\mem[24][12] ), .A2(n1149), .B1(\mem[26][12] ), .B2(
        n1148), .ZN(n929) );
  AOI22D0 U1786 ( .A1(\mem[25][12] ), .A2(n1151), .B1(\mem[27][12] ), .B2(
        n1150), .ZN(n928) );
  AOI22D0 U1787 ( .A1(\mem[21][12] ), .A2(n1159), .B1(\mem[23][12] ), .B2(
        n1158), .ZN(n934) );
  AOI22D0 U1788 ( .A1(\mem[28][12] ), .A2(n1161), .B1(\mem[30][12] ), .B2(
        n1160), .ZN(n933) );
  AOI22D0 U1789 ( .A1(\mem[29][12] ), .A2(n1163), .B1(\mem[31][12] ), .B2(
        n1162), .ZN(n932) );
  ND4D0 U1790 ( .A1(n935), .A2(n934), .A3(n933), .A4(n932), .ZN(n936) );
  OR4D0 U1791 ( .A1(n939), .A2(n938), .A3(n937), .A4(n936), .Z(A[12]) );
  AOI22D0 U1792 ( .A1(\mem[0][10] ), .A2(n1121), .B1(\mem[2][10] ), .B2(n1120), 
        .ZN(n943) );
  AOI22D0 U1793 ( .A1(\mem[1][10] ), .A2(n1123), .B1(\mem[3][10] ), .B2(n1122), 
        .ZN(n942) );
  AOI22D0 U1794 ( .A1(\mem[8][10] ), .A2(n1125), .B1(\mem[10][10] ), .B2(n1124), .ZN(n941) );
  AOI22D0 U1795 ( .A1(\mem[11][10] ), .A2(n1127), .B1(\mem[9][10] ), .B2(n1126), .ZN(n940) );
  ND4D0 U1796 ( .A1(n943), .A2(n942), .A3(n941), .A4(n940), .ZN(n959) );
  AOI22D0 U1797 ( .A1(\mem[4][10] ), .A2(n1133), .B1(\mem[6][10] ), .B2(n1132), 
        .ZN(n947) );
  AOI22D0 U1798 ( .A1(\mem[5][10] ), .A2(n1135), .B1(\mem[7][10] ), .B2(n1134), 
        .ZN(n946) );
  AOI22D0 U1799 ( .A1(\mem[12][10] ), .A2(n1137), .B1(\mem[14][10] ), .B2(
        n1136), .ZN(n945) );
  AOI22D0 U1800 ( .A1(\mem[13][10] ), .A2(n1139), .B1(\mem[15][10] ), .B2(
        n1138), .ZN(n944) );
  ND4D0 U1801 ( .A1(n947), .A2(n946), .A3(n945), .A4(n944), .ZN(n958) );
  AOI22D0 U1802 ( .A1(\mem[16][10] ), .A2(n1145), .B1(\mem[18][10] ), .B2(
        n1144), .ZN(n951) );
  AOI22D0 U1803 ( .A1(\mem[17][10] ), .A2(n1147), .B1(\mem[19][10] ), .B2(
        n1146), .ZN(n950) );
  AOI22D0 U1804 ( .A1(\mem[25][10] ), .A2(n1151), .B1(\mem[27][10] ), .B2(
        n1150), .ZN(n948) );
  ND4D0 U1805 ( .A1(n951), .A2(n950), .A3(n949), .A4(n948), .ZN(n957) );
  AOI22D0 U1806 ( .A1(\mem[20][10] ), .A2(n1157), .B1(\mem[22][10] ), .B2(
        n1156), .ZN(n955) );
  AOI22D0 U1807 ( .A1(\mem[21][10] ), .A2(n1159), .B1(\mem[23][10] ), .B2(
        n1158), .ZN(n954) );
  AOI22D0 U1808 ( .A1(\mem[28][10] ), .A2(n1161), .B1(\mem[30][10] ), .B2(
        n1160), .ZN(n953) );
  AOI22D0 U1809 ( .A1(\mem[29][10] ), .A2(n1163), .B1(\mem[31][10] ), .B2(
        n1162), .ZN(n952) );
  ND4D0 U1810 ( .A1(n955), .A2(n954), .A3(n953), .A4(n952), .ZN(n956) );
  OR4D0 U1811 ( .A1(n959), .A2(n958), .A3(n957), .A4(n956), .Z(A[10]) );
  AOI22D0 U1812 ( .A1(\mem[0][7] ), .A2(n1121), .B1(\mem[2][7] ), .B2(n1120), 
        .ZN(n963) );
  AOI22D0 U1813 ( .A1(\mem[1][7] ), .A2(n1123), .B1(\mem[3][7] ), .B2(n1122), 
        .ZN(n962) );
  AOI22D0 U1814 ( .A1(\mem[8][7] ), .A2(n1125), .B1(\mem[10][7] ), .B2(n1124), 
        .ZN(n961) );
  AOI22D0 U1815 ( .A1(\mem[11][7] ), .A2(n1127), .B1(\mem[9][7] ), .B2(n1126), 
        .ZN(n960) );
  ND4D0 U1816 ( .A1(n963), .A2(n962), .A3(n961), .A4(n960), .ZN(n979) );
  AOI22D0 U1817 ( .A1(\mem[4][7] ), .A2(n1133), .B1(\mem[6][7] ), .B2(n1132), 
        .ZN(n967) );
  AOI22D0 U1818 ( .A1(\mem[5][7] ), .A2(n1135), .B1(\mem[7][7] ), .B2(n1134), 
        .ZN(n966) );
  AOI22D0 U1819 ( .A1(\mem[12][7] ), .A2(n1137), .B1(\mem[14][7] ), .B2(n1136), 
        .ZN(n965) );
  ND4D0 U1820 ( .A1(n967), .A2(n966), .A3(n965), .A4(n964), .ZN(n978) );
  AOI22D0 U1821 ( .A1(\mem[16][7] ), .A2(n1145), .B1(\mem[18][7] ), .B2(n1144), 
        .ZN(n971) );
  AOI22D0 U1822 ( .A1(\mem[17][7] ), .A2(n1147), .B1(\mem[19][7] ), .B2(n1146), 
        .ZN(n970) );
  AOI22D0 U1823 ( .A1(\mem[24][7] ), .A2(n1149), .B1(\mem[26][7] ), .B2(n1148), 
        .ZN(n969) );
  AOI22D0 U1824 ( .A1(\mem[25][7] ), .A2(n1151), .B1(\mem[27][7] ), .B2(n1150), 
        .ZN(n968) );
  ND4D0 U1825 ( .A1(n971), .A2(n970), .A3(n969), .A4(n968), .ZN(n977) );
  AOI22D0 U1826 ( .A1(\mem[20][7] ), .A2(n1157), .B1(\mem[22][7] ), .B2(n1156), 
        .ZN(n975) );
  AOI22D0 U1827 ( .A1(\mem[21][7] ), .A2(n1159), .B1(\mem[23][7] ), .B2(n1158), 
        .ZN(n974) );
  AOI22D0 U1828 ( .A1(\mem[28][7] ), .A2(n1161), .B1(\mem[30][7] ), .B2(n1160), 
        .ZN(n973) );
  AOI22D0 U1829 ( .A1(\mem[29][7] ), .A2(n1163), .B1(\mem[31][7] ), .B2(n1162), 
        .ZN(n972) );
  ND4D0 U1830 ( .A1(n975), .A2(n974), .A3(n973), .A4(n972), .ZN(n976) );
  OR4D0 U1831 ( .A1(n979), .A2(n978), .A3(n977), .A4(n976), .Z(A[7]) );
  AOI22D0 U1832 ( .A1(\mem[0][6] ), .A2(n1121), .B1(\mem[2][6] ), .B2(n1120), 
        .ZN(n983) );
  AOI22D0 U1833 ( .A1(\mem[1][6] ), .A2(n1123), .B1(\mem[3][6] ), .B2(n1122), 
        .ZN(n982) );
  AOI22D0 U1834 ( .A1(\mem[8][6] ), .A2(n1125), .B1(\mem[10][6] ), .B2(n1124), 
        .ZN(n981) );
  AOI22D0 U1835 ( .A1(\mem[11][6] ), .A2(n1127), .B1(\mem[9][6] ), .B2(n1126), 
        .ZN(n980) );
  ND4D0 U1836 ( .A1(n983), .A2(n982), .A3(n981), .A4(n980), .ZN(n999) );
  AOI22D0 U1837 ( .A1(\mem[4][6] ), .A2(n1133), .B1(\mem[6][6] ), .B2(n1132), 
        .ZN(n987) );
  AOI22D0 U1838 ( .A1(\mem[5][6] ), .A2(n1135), .B1(\mem[7][6] ), .B2(n1134), 
        .ZN(n986) );
  AOI22D0 U1839 ( .A1(\mem[13][6] ), .A2(n1139), .B1(\mem[15][6] ), .B2(n1138), 
        .ZN(n984) );
  ND4D0 U1840 ( .A1(n987), .A2(n986), .A3(n985), .A4(n984), .ZN(n998) );
  AOI22D0 U1841 ( .A1(\mem[16][6] ), .A2(n1145), .B1(\mem[18][6] ), .B2(n1144), 
        .ZN(n991) );
  AOI22D0 U1842 ( .A1(\mem[17][6] ), .A2(n1147), .B1(\mem[19][6] ), .B2(n1146), 
        .ZN(n990) );
  AOI22D0 U1843 ( .A1(\mem[24][6] ), .A2(n1149), .B1(\mem[26][6] ), .B2(n1148), 
        .ZN(n989) );
  AOI22D0 U1844 ( .A1(\mem[25][6] ), .A2(n1151), .B1(\mem[27][6] ), .B2(n1150), 
        .ZN(n988) );
  ND4D0 U1845 ( .A1(n991), .A2(n990), .A3(n989), .A4(n988), .ZN(n997) );
  AOI22D0 U1846 ( .A1(\mem[20][6] ), .A2(n1157), .B1(\mem[22][6] ), .B2(n1156), 
        .ZN(n995) );
  AOI22D0 U1847 ( .A1(\mem[21][6] ), .A2(n1159), .B1(\mem[23][6] ), .B2(n1158), 
        .ZN(n994) );
  AOI22D0 U1848 ( .A1(\mem[28][6] ), .A2(n1161), .B1(\mem[30][6] ), .B2(n1160), 
        .ZN(n993) );
  AOI22D0 U1849 ( .A1(\mem[29][6] ), .A2(n1163), .B1(\mem[31][6] ), .B2(n1162), 
        .ZN(n992) );
  ND4D0 U1850 ( .A1(n995), .A2(n994), .A3(n993), .A4(n992), .ZN(n996) );
  OR4D0 U1851 ( .A1(n999), .A2(n998), .A3(n997), .A4(n996), .Z(A[6]) );
  AOI22D0 U1852 ( .A1(\mem[0][4] ), .A2(n1121), .B1(\mem[2][4] ), .B2(n1120), 
        .ZN(n1003) );
  AOI22D0 U1853 ( .A1(\mem[1][4] ), .A2(n1123), .B1(\mem[3][4] ), .B2(n1122), 
        .ZN(n1002) );
  AOI22D0 U1854 ( .A1(\mem[8][4] ), .A2(n1125), .B1(\mem[10][4] ), .B2(n1124), 
        .ZN(n1001) );
  AOI22D0 U1855 ( .A1(\mem[11][4] ), .A2(n1127), .B1(\mem[9][4] ), .B2(n1126), 
        .ZN(n1000) );
  AOI22D0 U1856 ( .A1(\mem[5][4] ), .A2(n1135), .B1(\mem[7][4] ), .B2(n1134), 
        .ZN(n1006) );
  AOI22D0 U1857 ( .A1(\mem[12][4] ), .A2(n1137), .B1(\mem[14][4] ), .B2(n1136), 
        .ZN(n1005) );
  AOI22D0 U1858 ( .A1(\mem[13][4] ), .A2(n1139), .B1(\mem[15][4] ), .B2(n1138), 
        .ZN(n1004) );
  ND4D0 U1859 ( .A1(n1007), .A2(n1006), .A3(n1005), .A4(n1004), .ZN(n1018) );
  AOI22D0 U1860 ( .A1(\mem[16][4] ), .A2(n1145), .B1(\mem[18][4] ), .B2(n1144), 
        .ZN(n1011) );
  AOI22D0 U1861 ( .A1(\mem[17][4] ), .A2(n1147), .B1(\mem[19][4] ), .B2(n1146), 
        .ZN(n1010) );
  AOI22D0 U1862 ( .A1(\mem[24][4] ), .A2(n1149), .B1(\mem[26][4] ), .B2(n1148), 
        .ZN(n1009) );
  AOI22D0 U1863 ( .A1(\mem[25][4] ), .A2(n1151), .B1(\mem[27][4] ), .B2(n1150), 
        .ZN(n1008) );
  ND4D0 U1864 ( .A1(n1011), .A2(n1010), .A3(n1009), .A4(n1008), .ZN(n1017) );
  AOI22D0 U1865 ( .A1(\mem[20][4] ), .A2(n1157), .B1(\mem[22][4] ), .B2(n1156), 
        .ZN(n1015) );
  AOI22D0 U1866 ( .A1(\mem[21][4] ), .A2(n1159), .B1(\mem[23][4] ), .B2(n1158), 
        .ZN(n1014) );
  AOI22D0 U1867 ( .A1(\mem[28][4] ), .A2(n1161), .B1(\mem[30][4] ), .B2(n1160), 
        .ZN(n1013) );
  AOI22D0 U1868 ( .A1(\mem[29][4] ), .A2(n1163), .B1(\mem[31][4] ), .B2(n1162), 
        .ZN(n1012) );
  ND4D0 U1869 ( .A1(n1015), .A2(n1014), .A3(n1013), .A4(n1012), .ZN(n1016) );
  OR4D0 U1870 ( .A1(n1019), .A2(n1018), .A3(n1017), .A4(n1016), .Z(A[4]) );
  AOI22D0 U1871 ( .A1(\mem[0][1] ), .A2(n1121), .B1(\mem[2][1] ), .B2(n1120), 
        .ZN(n1023) );
  AOI22D0 U1872 ( .A1(\mem[8][1] ), .A2(n1125), .B1(\mem[10][1] ), .B2(n1124), 
        .ZN(n1021) );
  AOI22D0 U1873 ( .A1(\mem[11][1] ), .A2(n1127), .B1(\mem[9][1] ), .B2(n1126), 
        .ZN(n1020) );
  ND4D0 U1874 ( .A1(n1023), .A2(n1022), .A3(n1021), .A4(n1020), .ZN(n1039) );
  AOI22D0 U1875 ( .A1(\mem[4][1] ), .A2(n1133), .B1(\mem[6][1] ), .B2(n1132), 
        .ZN(n1027) );
  AOI22D0 U1876 ( .A1(\mem[5][1] ), .A2(n1135), .B1(\mem[7][1] ), .B2(n1134), 
        .ZN(n1026) );
  AOI22D0 U1877 ( .A1(\mem[12][1] ), .A2(n1137), .B1(\mem[14][1] ), .B2(n1136), 
        .ZN(n1025) );
  AOI22D0 U1878 ( .A1(\mem[13][1] ), .A2(n1139), .B1(\mem[15][1] ), .B2(n1138), 
        .ZN(n1024) );
  ND4D0 U1879 ( .A1(n1027), .A2(n1026), .A3(n1025), .A4(n1024), .ZN(n1038) );
  AOI22D0 U1880 ( .A1(\mem[16][1] ), .A2(n1145), .B1(\mem[18][1] ), .B2(n1144), 
        .ZN(n1031) );
  AOI22D0 U1881 ( .A1(\mem[17][1] ), .A2(n1147), .B1(\mem[19][1] ), .B2(n1146), 
        .ZN(n1030) );
  AOI22D0 U1882 ( .A1(\mem[24][1] ), .A2(n1149), .B1(\mem[26][1] ), .B2(n1148), 
        .ZN(n1029) );
  AOI22D0 U1883 ( .A1(\mem[25][1] ), .A2(n1151), .B1(\mem[27][1] ), .B2(n1150), 
        .ZN(n1028) );
  ND4D0 U1884 ( .A1(n1031), .A2(n1030), .A3(n1029), .A4(n1028), .ZN(n1037) );
  AOI22D0 U1885 ( .A1(\mem[20][1] ), .A2(n1157), .B1(\mem[22][1] ), .B2(n1156), 
        .ZN(n1035) );
  AOI22D0 U1886 ( .A1(\mem[21][1] ), .A2(n1159), .B1(\mem[23][1] ), .B2(n1158), 
        .ZN(n1034) );
  AOI22D0 U1887 ( .A1(\mem[28][1] ), .A2(n1161), .B1(\mem[30][1] ), .B2(n1160), 
        .ZN(n1033) );
  AOI22D0 U1888 ( .A1(\mem[29][1] ), .A2(n1163), .B1(\mem[31][1] ), .B2(n1162), 
        .ZN(n1032) );
  OR4D0 U1889 ( .A1(n1039), .A2(n1038), .A3(n1037), .A4(n1036), .Z(A[1]) );
  AOI22D0 U1890 ( .A1(\mem[0][0] ), .A2(n1121), .B1(\mem[2][0] ), .B2(n1120), 
        .ZN(n1043) );
  AOI22D0 U1891 ( .A1(\mem[1][0] ), .A2(n1123), .B1(\mem[3][0] ), .B2(n1122), 
        .ZN(n1042) );
  AOI22D0 U1892 ( .A1(\mem[8][0] ), .A2(n1125), .B1(\mem[10][0] ), .B2(n1124), 
        .ZN(n1041) );
  AOI22D0 U1893 ( .A1(\mem[11][0] ), .A2(n1127), .B1(\mem[9][0] ), .B2(n1126), 
        .ZN(n1040) );
  ND4D0 U1894 ( .A1(n1043), .A2(n1042), .A3(n1041), .A4(n1040), .ZN(n1059) );
  AOI22D0 U1895 ( .A1(\mem[4][0] ), .A2(n1133), .B1(\mem[6][0] ), .B2(n1132), 
        .ZN(n1047) );
  AOI22D0 U1896 ( .A1(\mem[12][0] ), .A2(n1137), .B1(\mem[14][0] ), .B2(n1136), 
        .ZN(n1045) );
  AOI22D0 U1897 ( .A1(\mem[13][0] ), .A2(n1139), .B1(\mem[15][0] ), .B2(n1138), 
        .ZN(n1044) );
  ND4D0 U1898 ( .A1(n1047), .A2(n1046), .A3(n1045), .A4(n1044), .ZN(n1058) );
  AOI22D0 U1899 ( .A1(\mem[16][0] ), .A2(n1145), .B1(\mem[18][0] ), .B2(n1144), 
        .ZN(n1051) );
  AOI22D0 U1900 ( .A1(\mem[17][0] ), .A2(n1147), .B1(\mem[19][0] ), .B2(n1146), 
        .ZN(n1050) );
  AOI22D0 U1901 ( .A1(\mem[24][0] ), .A2(n1149), .B1(\mem[26][0] ), .B2(n1148), 
        .ZN(n1049) );
  AOI22D0 U1902 ( .A1(\mem[25][0] ), .A2(n1151), .B1(\mem[27][0] ), .B2(n1150), 
        .ZN(n1048) );
  ND4D0 U1903 ( .A1(n1051), .A2(n1050), .A3(n1049), .A4(n1048), .ZN(n1057) );
  AOI22D0 U1904 ( .A1(\mem[20][0] ), .A2(n1157), .B1(\mem[22][0] ), .B2(n1156), 
        .ZN(n1055) );
  AOI22D0 U1905 ( .A1(\mem[21][0] ), .A2(n1159), .B1(\mem[23][0] ), .B2(n1158), 
        .ZN(n1054) );
  AOI22D0 U1906 ( .A1(\mem[28][0] ), .A2(n1161), .B1(\mem[30][0] ), .B2(n1160), 
        .ZN(n1053) );
  AOI22D0 U1907 ( .A1(\mem[29][0] ), .A2(n1163), .B1(\mem[31][0] ), .B2(n1162), 
        .ZN(n1052) );
  ND4D0 U1908 ( .A1(n1055), .A2(n1054), .A3(n1053), .A4(n1052), .ZN(n1056) );
  OR4D0 U1909 ( .A1(n1059), .A2(n1058), .A3(n1057), .A4(n1056), .Z(A[0]) );
  AOI22D0 U1910 ( .A1(\mem[0][3] ), .A2(n1121), .B1(\mem[2][3] ), .B2(n1120), 
        .ZN(n1063) );
  AOI22D0 U1911 ( .A1(\mem[1][3] ), .A2(n1123), .B1(\mem[3][3] ), .B2(n1122), 
        .ZN(n1062) );
  AOI22D0 U1912 ( .A1(\mem[8][3] ), .A2(n1125), .B1(\mem[10][3] ), .B2(n1124), 
        .ZN(n1061) );
  ND4D0 U1913 ( .A1(n1063), .A2(n1062), .A3(n1061), .A4(n1060), .ZN(n1079) );
  AOI22D0 U1914 ( .A1(\mem[4][3] ), .A2(n1133), .B1(\mem[6][3] ), .B2(n1132), 
        .ZN(n1067) );
  AOI22D0 U1915 ( .A1(\mem[5][3] ), .A2(n1135), .B1(\mem[7][3] ), .B2(n1134), 
        .ZN(n1066) );
  AOI22D0 U1916 ( .A1(\mem[12][3] ), .A2(n1137), .B1(\mem[14][3] ), .B2(n1136), 
        .ZN(n1065) );
  AOI22D0 U1917 ( .A1(\mem[13][3] ), .A2(n1139), .B1(\mem[15][3] ), .B2(n1138), 
        .ZN(n1064) );
  ND4D0 U1918 ( .A1(n1067), .A2(n1066), .A3(n1065), .A4(n1064), .ZN(n1078) );
  AOI22D0 U1919 ( .A1(\mem[16][3] ), .A2(n1145), .B1(\mem[18][3] ), .B2(n1144), 
        .ZN(n1071) );
  AOI22D0 U1920 ( .A1(\mem[17][3] ), .A2(n1147), .B1(\mem[19][3] ), .B2(n1146), 
        .ZN(n1070) );
  AOI22D0 U1921 ( .A1(\mem[24][3] ), .A2(n1149), .B1(\mem[26][3] ), .B2(n1148), 
        .ZN(n1069) );
  AOI22D0 U1922 ( .A1(\mem[25][3] ), .A2(n1151), .B1(\mem[27][3] ), .B2(n1150), 
        .ZN(n1068) );
  ND4D0 U1923 ( .A1(n1071), .A2(n1070), .A3(n1069), .A4(n1068), .ZN(n1077) );
  AOI22D0 U1924 ( .A1(\mem[20][3] ), .A2(n1157), .B1(\mem[22][3] ), .B2(n1156), 
        .ZN(n1075) );
  AOI22D0 U1925 ( .A1(\mem[21][3] ), .A2(n1159), .B1(\mem[23][3] ), .B2(n1158), 
        .ZN(n1074) );
  AOI22D0 U1926 ( .A1(\mem[28][3] ), .A2(n1161), .B1(\mem[30][3] ), .B2(n1160), 
        .ZN(n1073) );
  AOI22D0 U1927 ( .A1(\mem[29][3] ), .A2(n1163), .B1(\mem[31][3] ), .B2(n1162), 
        .ZN(n1072) );
  ND4D0 U1928 ( .A1(n1075), .A2(n1074), .A3(n1073), .A4(n1072), .ZN(n1076) );
  OR4D0 U1929 ( .A1(n1079), .A2(n1078), .A3(n1077), .A4(n1076), .Z(A[3]) );
  AOI22D0 U1930 ( .A1(\mem[0][9] ), .A2(n1121), .B1(\mem[2][9] ), .B2(n1120), 
        .ZN(n1083) );
  AOI22D0 U1931 ( .A1(\mem[1][9] ), .A2(n1123), .B1(\mem[3][9] ), .B2(n1122), 
        .ZN(n1082) );
  AOI22D0 U1932 ( .A1(\mem[8][9] ), .A2(n1125), .B1(\mem[10][9] ), .B2(n1124), 
        .ZN(n1081) );
  AOI22D0 U1933 ( .A1(\mem[11][9] ), .A2(n1127), .B1(\mem[9][9] ), .B2(n1126), 
        .ZN(n1080) );
  ND4D0 U1934 ( .A1(n1083), .A2(n1082), .A3(n1081), .A4(n1080), .ZN(n1099) );
  AOI22D0 U1935 ( .A1(\mem[4][9] ), .A2(n1133), .B1(\mem[6][9] ), .B2(n1132), 
        .ZN(n1087) );
  AOI22D0 U1936 ( .A1(\mem[5][9] ), .A2(n1135), .B1(\mem[7][9] ), .B2(n1134), 
        .ZN(n1086) );
  AOI22D0 U1937 ( .A1(\mem[12][9] ), .A2(n1137), .B1(\mem[14][9] ), .B2(n1136), 
        .ZN(n1085) );
  AOI22D0 U1938 ( .A1(\mem[13][9] ), .A2(n1139), .B1(\mem[15][9] ), .B2(n1138), 
        .ZN(n1084) );
  ND4D0 U1939 ( .A1(n1087), .A2(n1086), .A3(n1085), .A4(n1084), .ZN(n1098) );
  AOI22D0 U1940 ( .A1(\mem[16][9] ), .A2(n1145), .B1(\mem[18][9] ), .B2(n1144), 
        .ZN(n1091) );
  AOI22D0 U1941 ( .A1(\mem[24][9] ), .A2(n1149), .B1(\mem[26][9] ), .B2(n1148), 
        .ZN(n1089) );
  AOI22D0 U1942 ( .A1(\mem[25][9] ), .A2(n1151), .B1(\mem[27][9] ), .B2(n1150), 
        .ZN(n1088) );
  ND4D0 U1943 ( .A1(n1091), .A2(n1090), .A3(n1089), .A4(n1088), .ZN(n1097) );
  AOI22D0 U1944 ( .A1(\mem[20][9] ), .A2(n1157), .B1(\mem[22][9] ), .B2(n1156), 
        .ZN(n1095) );
  AOI22D0 U1945 ( .A1(\mem[21][9] ), .A2(n1159), .B1(\mem[23][9] ), .B2(n1158), 
        .ZN(n1094) );
  AOI22D0 U1946 ( .A1(\mem[28][9] ), .A2(n1161), .B1(\mem[30][9] ), .B2(n1160), 
        .ZN(n1093) );
  AOI22D0 U1947 ( .A1(\mem[29][9] ), .A2(n1163), .B1(\mem[31][9] ), .B2(n1162), 
        .ZN(n1092) );
  ND4D0 U1948 ( .A1(n1095), .A2(n1094), .A3(n1093), .A4(n1092), .ZN(n1096) );
  OR4D0 U1949 ( .A1(n1099), .A2(n1098), .A3(n1097), .A4(n1096), .Z(A[9]) );
  AOI22D0 U1950 ( .A1(\mem[1][15] ), .A2(n1123), .B1(\mem[3][15] ), .B2(n1122), 
        .ZN(n1102) );
  AOI22D0 U1951 ( .A1(\mem[8][15] ), .A2(n1125), .B1(\mem[10][15] ), .B2(n1124), .ZN(n1101) );
  AOI22D0 U1952 ( .A1(\mem[11][15] ), .A2(n1127), .B1(\mem[9][15] ), .B2(n1126), .ZN(n1100) );
  ND4D0 U1953 ( .A1(n1103), .A2(n1102), .A3(n1101), .A4(n1100), .ZN(n1119) );
  AOI22D0 U1954 ( .A1(\mem[4][15] ), .A2(n1133), .B1(\mem[6][15] ), .B2(n1132), 
        .ZN(n1107) );
  AOI22D0 U1955 ( .A1(\mem[5][15] ), .A2(n1135), .B1(\mem[7][15] ), .B2(n1134), 
        .ZN(n1106) );
  AOI22D0 U1956 ( .A1(\mem[12][15] ), .A2(n1137), .B1(\mem[14][15] ), .B2(
        n1136), .ZN(n1105) );
  AOI22D0 U1957 ( .A1(\mem[13][15] ), .A2(n1139), .B1(\mem[15][15] ), .B2(
        n1138), .ZN(n1104) );
  ND4D0 U1958 ( .A1(n1107), .A2(n1106), .A3(n1105), .A4(n1104), .ZN(n1118) );
  AOI22D0 U1959 ( .A1(\mem[16][15] ), .A2(n1145), .B1(\mem[18][15] ), .B2(
        n1144), .ZN(n1111) );
  AOI22D0 U1960 ( .A1(\mem[17][15] ), .A2(n1147), .B1(\mem[19][15] ), .B2(
        n1146), .ZN(n1110) );
  AOI22D0 U1961 ( .A1(\mem[24][15] ), .A2(n1149), .B1(\mem[26][15] ), .B2(
        n1148), .ZN(n1109) );
  AOI22D0 U1962 ( .A1(\mem[25][15] ), .A2(n1151), .B1(\mem[27][15] ), .B2(
        n1150), .ZN(n1108) );
  ND4D0 U1963 ( .A1(n1111), .A2(n1110), .A3(n1109), .A4(n1108), .ZN(n1117) );
  AOI22D0 U1964 ( .A1(\mem[20][15] ), .A2(n1157), .B1(\mem[22][15] ), .B2(
        n1156), .ZN(n1115) );
  AOI22D0 U1965 ( .A1(\mem[21][15] ), .A2(n1159), .B1(\mem[23][15] ), .B2(
        n1158), .ZN(n1114) );
  AOI22D0 U1966 ( .A1(\mem[28][15] ), .A2(n1161), .B1(\mem[30][15] ), .B2(
        n1160), .ZN(n1113) );
  ND4D0 U1967 ( .A1(n1115), .A2(n1114), .A3(n1113), .A4(n1112), .ZN(n1116) );
  OR4D0 U1968 ( .A1(n1119), .A2(n1118), .A3(n1117), .A4(n1116), .Z(A[15]) );
  AOI22D0 U1969 ( .A1(\mem[0][21] ), .A2(n1121), .B1(\mem[2][21] ), .B2(n1120), 
        .ZN(n1131) );
  AOI22D0 U1970 ( .A1(\mem[1][21] ), .A2(n1123), .B1(\mem[3][21] ), .B2(n1122), 
        .ZN(n1130) );
  AOI22D0 U1971 ( .A1(\mem[8][21] ), .A2(n1125), .B1(\mem[10][21] ), .B2(n1124), .ZN(n1129) );
  AOI22D0 U1972 ( .A1(\mem[11][21] ), .A2(n1127), .B1(\mem[9][21] ), .B2(n1126), .ZN(n1128) );
  ND4D0 U1973 ( .A1(n1131), .A2(n1130), .A3(n1129), .A4(n1128), .ZN(n1939) );
  AOI22D0 U1974 ( .A1(\mem[4][21] ), .A2(n1133), .B1(\mem[6][21] ), .B2(n1132), 
        .ZN(n1143) );
  AOI22D0 U1975 ( .A1(\mem[5][21] ), .A2(n1135), .B1(\mem[7][21] ), .B2(n1134), 
        .ZN(n1142) );
  AOI22D0 U1976 ( .A1(\mem[13][21] ), .A2(n1139), .B1(\mem[15][21] ), .B2(
        n1138), .ZN(n1140) );
  ND4D0 U1977 ( .A1(n1143), .A2(n1142), .A3(n1141), .A4(n1140), .ZN(n1938) );
  AOI22D0 U1978 ( .A1(\mem[16][21] ), .A2(n1145), .B1(\mem[18][21] ), .B2(
        n1144), .ZN(n1155) );
  AOI22D0 U1979 ( .A1(\mem[17][21] ), .A2(n1147), .B1(\mem[19][21] ), .B2(
        n1146), .ZN(n1154) );
  AOI22D0 U1980 ( .A1(\mem[24][21] ), .A2(n1149), .B1(\mem[26][21] ), .B2(
        n1148), .ZN(n1153) );
  AOI22D0 U1981 ( .A1(\mem[25][21] ), .A2(n1151), .B1(\mem[27][21] ), .B2(
        n1150), .ZN(n1152) );
  ND4D0 U1982 ( .A1(n1155), .A2(n1154), .A3(n1153), .A4(n1152), .ZN(n1169) );
  AOI22D0 U1983 ( .A1(\mem[20][21] ), .A2(n1157), .B1(\mem[22][21] ), .B2(
        n1156), .ZN(n1167) );
  AOI22D0 U1984 ( .A1(\mem[21][21] ), .A2(n1159), .B1(\mem[23][21] ), .B2(
        n1158), .ZN(n1166) );
  AOI22D0 U1985 ( .A1(\mem[28][21] ), .A2(n1161), .B1(\mem[30][21] ), .B2(
        n1160), .ZN(n1165) );
  AOI22D0 U1986 ( .A1(\mem[29][21] ), .A2(n1163), .B1(\mem[31][21] ), .B2(
        n1162), .ZN(n1164) );
  ND4D0 U1987 ( .A1(n1167), .A2(n1166), .A3(n1165), .A4(n1164), .ZN(n1168) );
  OR4D0 U1988 ( .A1(n1939), .A2(n1938), .A3(n1169), .A4(n1168), .Z(A[21]) );
endmodule
