// Created by ihdl
module rom_256x16 ( clk, addr, dout, prog_we, prog_addr, prog_data );
  input [7:0] addr;
  output [15:0] dout;
  input [7:0] prog_addr;
  input [15:0] prog_data;
  input clk, prog_we;
  wire   \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , \mem[1][15] , \mem[1][14] , \mem[1][13] , \mem[1][12] ,
         \mem[1][11] , \mem[1][10] , \mem[1][9] , \mem[1][8] , \mem[1][7] ,
         \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] ,
         \mem[1][1] , \mem[1][0] , \mem[2][15] , \mem[2][14] , \mem[2][13] ,
         \mem[2][12] , \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] ,
         \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] ,
         \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[3][15] , \mem[3][14] ,
         \mem[3][13] , \mem[3][12] , \mem[3][11] , \mem[3][10] , \mem[3][9] ,
         \mem[3][8] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[4][15] ,
         \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] , \mem[4][10] ,
         \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] , \mem[4][5] ,
         \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] , \mem[4][0] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[6][15] , \mem[6][14] , \mem[6][13] , \mem[6][12] ,
         \mem[6][11] , \mem[6][10] , \mem[6][9] , \mem[6][8] , \mem[6][7] ,
         \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] ,
         \mem[6][1] , \mem[6][0] , \mem[7][15] , \mem[7][14] , \mem[7][13] ,
         \mem[7][12] , \mem[7][11] , \mem[7][10] , \mem[7][9] , \mem[7][8] ,
         \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] ,
         \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[8][15] , \mem[8][14] ,
         \mem[8][13] , \mem[8][12] , \mem[8][11] , \mem[8][10] , \mem[8][9] ,
         \mem[8][8] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[9][15] ,
         \mem[9][14] , \mem[9][13] , \mem[9][12] , \mem[9][11] , \mem[9][10] ,
         \mem[9][9] , \mem[9][8] , \mem[9][7] , \mem[9][6] , \mem[9][5] ,
         \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] , \mem[9][0] ,
         \mem[10][15] , \mem[10][14] , \mem[10][13] , \mem[10][12] ,
         \mem[10][11] , \mem[10][10] , \mem[10][9] , \mem[10][8] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[11][15] ,
         \mem[11][14] , \mem[11][13] , \mem[11][12] , \mem[11][11] ,
         \mem[11][10] , \mem[11][9] , \mem[11][8] , \mem[11][7] , \mem[11][6] ,
         \mem[11][5] , \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] ,
         \mem[11][0] , \mem[12][15] , \mem[12][14] , \mem[12][13] ,
         \mem[12][12] , \mem[12][11] , \mem[12][10] , \mem[12][9] ,
         \mem[12][8] , \mem[12][7] , \mem[12][6] , \mem[12][5] , \mem[12][4] ,
         \mem[12][3] , \mem[12][2] , \mem[12][1] , \mem[12][0] , \mem[13][15] ,
         \mem[13][14] , \mem[13][13] , \mem[13][12] , \mem[13][11] ,
         \mem[13][10] , \mem[13][9] , \mem[13][8] , \mem[13][7] , \mem[13][6] ,
         \mem[13][5] , \mem[13][4] , \mem[13][3] , \mem[13][2] , \mem[13][1] ,
         \mem[13][0] , \mem[14][15] , \mem[14][14] , \mem[14][13] ,
         \mem[14][12] , \mem[14][11] , \mem[14][10] , \mem[14][9] ,
         \mem[14][8] , \mem[14][7] , \mem[14][6] , \mem[14][5] , \mem[14][4] ,
         \mem[14][3] , \mem[14][2] , \mem[14][1] , \mem[14][0] , \mem[15][15] ,
         \mem[15][14] , \mem[15][13] , \mem[15][12] , \mem[15][11] ,
         \mem[15][10] , \mem[15][9] , \mem[15][8] , \mem[15][7] , \mem[15][6] ,
         \mem[15][5] , \mem[15][4] , \mem[15][3] , \mem[15][2] , \mem[15][1] ,
         \mem[15][0] , \mem[16][15] , \mem[16][14] , \mem[16][13] ,
         \mem[16][12] , \mem[16][11] , \mem[16][10] , \mem[16][9] ,
         \mem[16][8] , \mem[16][7] , \mem[16][6] , \mem[16][5] , \mem[16][4] ,
         \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] , \mem[17][15] ,
         \mem[17][14] , \mem[17][13] , \mem[17][12] , \mem[17][11] ,
         \mem[17][10] , \mem[17][9] , \mem[17][8] , \mem[17][7] , \mem[17][6] ,
         \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] , \mem[17][1] ,
         \mem[17][0] , \mem[18][15] , \mem[18][14] , \mem[18][13] ,
         \mem[18][12] , \mem[18][11] , \mem[18][10] , \mem[18][9] ,
         \mem[18][8] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[19][15] ,
         \mem[19][14] , \mem[19][13] , \mem[19][12] , \mem[19][11] ,
         \mem[19][10] , \mem[19][9] , \mem[19][8] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[20][15] , \mem[20][14] , \mem[20][13] ,
         \mem[20][12] , \mem[20][11] , \mem[20][10] , \mem[20][9] ,
         \mem[20][8] , \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] ,
         \mem[20][3] , \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[21][15] ,
         \mem[21][14] , \mem[21][13] , \mem[21][12] , \mem[21][11] ,
         \mem[21][10] , \mem[21][9] , \mem[21][8] , \mem[21][7] , \mem[21][6] ,
         \mem[21][5] , \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] ,
         \mem[21][0] , \mem[22][15] , \mem[22][14] , \mem[22][13] ,
         \mem[22][12] , \mem[22][11] , \mem[22][10] , \mem[22][9] ,
         \mem[22][8] , \mem[22][7] , \mem[22][6] , \mem[22][5] , \mem[22][4] ,
         \mem[22][3] , \mem[22][2] , \mem[22][1] , \mem[22][0] , \mem[23][15] ,
         \mem[23][14] , \mem[23][13] , \mem[23][12] , \mem[23][11] ,
         \mem[23][10] , \mem[23][9] , \mem[23][8] , \mem[23][7] , \mem[23][6] ,
         \mem[23][5] , \mem[23][4] , \mem[23][3] , \mem[23][2] , \mem[23][1] ,
         \mem[23][0] , \mem[24][15] , \mem[24][14] , \mem[24][13] ,
         \mem[24][12] , \mem[24][11] , \mem[24][10] , \mem[24][9] ,
         \mem[24][8] , \mem[24][7] , \mem[24][6] , \mem[24][5] , \mem[24][4] ,
         \mem[24][3] , \mem[24][2] , \mem[24][1] , \mem[24][0] , \mem[25][15] ,
         \mem[25][14] , \mem[25][13] , \mem[25][12] , \mem[25][11] ,
         \mem[25][10] , \mem[25][9] , \mem[25][8] , \mem[25][7] , \mem[25][6] ,
         \mem[25][5] , \mem[25][4] , \mem[25][3] , \mem[25][2] , \mem[25][1] ,
         \mem[25][0] , \mem[26][15] , \mem[26][14] , \mem[26][13] ,
         \mem[26][12] , \mem[26][11] , \mem[26][10] , \mem[26][9] ,
         \mem[26][8] , \mem[26][7] , \mem[26][6] , \mem[26][5] , \mem[26][4] ,
         \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] , \mem[27][15] ,
         \mem[27][14] , \mem[27][13] , \mem[27][12] , \mem[27][11] ,
         \mem[27][10] , \mem[27][9] , \mem[27][8] , \mem[27][7] , \mem[27][6] ,
         \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] , \mem[27][1] ,
         \mem[27][0] , \mem[28][15] , \mem[28][14] , \mem[28][13] ,
         \mem[28][12] , \mem[28][11] , \mem[28][10] , \mem[28][9] ,
         \mem[28][8] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[29][15] ,
         \mem[29][14] , \mem[29][13] , \mem[29][12] , \mem[29][11] ,
         \mem[29][10] , \mem[29][9] , \mem[29][8] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[30][15] , \mem[30][14] , \mem[30][13] ,
         \mem[30][12] , \mem[30][11] , \mem[30][10] , \mem[30][9] ,
         \mem[30][8] , \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] ,
         \mem[30][3] , \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[31][15] ,
         \mem[31][14] , \mem[31][13] , \mem[31][12] , \mem[31][11] ,
         \mem[31][10] , \mem[31][9] , \mem[31][8] , \mem[31][7] , \mem[31][6] ,
         \mem[31][5] , \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] ,
         \mem[31][0] , \mem[32][15] , \mem[32][14] , \mem[32][13] ,
         \mem[32][12] , \mem[32][11] , \mem[32][10] , \mem[32][9] ,
         \mem[32][8] , \mem[32][7] , \mem[32][6] , \mem[32][5] , \mem[32][4] ,
         \mem[32][3] , \mem[32][2] , \mem[32][1] , \mem[32][0] , \mem[33][15] ,
         \mem[33][14] , \mem[33][13] , \mem[33][12] , \mem[33][11] ,
         \mem[33][10] , \mem[33][9] , \mem[33][8] , \mem[33][7] , \mem[33][6] ,
         \mem[33][5] , \mem[33][4] , \mem[33][3] , \mem[33][2] , \mem[33][1] ,
         \mem[33][0] , \mem[34][15] , \mem[34][14] , \mem[34][13] ,
         \mem[34][12] , \mem[34][11] , \mem[34][10] , \mem[34][9] ,
         \mem[34][8] , \mem[34][7] , \mem[34][6] , \mem[34][5] , \mem[34][4] ,
         \mem[34][3] , \mem[34][2] , \mem[34][1] , \mem[34][0] , \mem[35][15] ,
         \mem[35][14] , \mem[35][13] , \mem[35][12] , \mem[35][11] ,
         \mem[35][10] , \mem[35][9] , \mem[35][8] , \mem[35][7] , \mem[35][6] ,
         \mem[35][5] , \mem[35][4] , \mem[35][3] , \mem[35][2] , \mem[35][1] ,
         \mem[35][0] , \mem[36][15] , \mem[36][14] , \mem[36][13] ,
         \mem[36][12] , \mem[36][11] , \mem[36][10] , \mem[36][9] ,
         \mem[36][8] , \mem[36][7] , \mem[36][6] , \mem[36][5] , \mem[36][4] ,
         \mem[36][3] , \mem[36][2] , \mem[36][1] , \mem[36][0] , \mem[37][15] ,
         \mem[37][14] , \mem[37][13] , \mem[37][12] , \mem[37][11] ,
         \mem[37][10] , \mem[37][9] , \mem[37][8] , \mem[37][7] , \mem[37][6] ,
         \mem[37][5] , \mem[37][4] , \mem[37][3] , \mem[37][2] , \mem[37][1] ,
         \mem[37][0] , \mem[38][15] , \mem[38][14] , \mem[38][13] ,
         \mem[38][12] , \mem[38][11] , \mem[38][10] , \mem[38][9] ,
         \mem[38][8] , \mem[38][7] , \mem[38][6] , \mem[38][5] , \mem[38][4] ,
         \mem[38][3] , \mem[38][2] , \mem[38][1] , \mem[38][0] , \mem[39][15] ,
         \mem[39][14] , \mem[39][13] , \mem[39][12] , \mem[39][11] ,
         \mem[39][10] , \mem[39][9] , \mem[39][8] , \mem[39][7] , \mem[39][6] ,
         \mem[39][5] , \mem[39][4] , \mem[39][3] , \mem[39][2] , \mem[39][1] ,
         \mem[39][0] , \mem[40][15] , \mem[40][14] , \mem[40][13] ,
         \mem[40][12] , \mem[40][11] , \mem[40][10] , \mem[40][9] ,
         \mem[40][8] , \mem[40][7] , \mem[40][6] , \mem[40][5] , \mem[40][4] ,
         \mem[40][3] , \mem[40][2] , \mem[40][1] , \mem[40][0] , \mem[41][15] ,
         \mem[41][14] , \mem[41][13] , \mem[41][12] , \mem[41][11] ,
         \mem[41][10] , \mem[41][9] , \mem[41][8] , \mem[41][7] , \mem[41][6] ,
         \mem[41][5] , \mem[41][4] , \mem[41][3] , \mem[41][2] , \mem[41][1] ,
         \mem[41][0] , \mem[42][15] , \mem[42][14] , \mem[42][13] ,
         \mem[42][12] , \mem[42][11] , \mem[42][10] , \mem[42][9] ,
         \mem[42][8] , \mem[42][7] , \mem[42][6] , \mem[42][5] , \mem[42][4] ,
         \mem[42][3] , \mem[42][2] , \mem[42][1] , \mem[42][0] , \mem[43][15] ,
         \mem[43][14] , \mem[43][13] , \mem[43][12] , \mem[43][11] ,
         \mem[43][10] , \mem[43][9] , \mem[43][8] , \mem[43][7] , \mem[43][6] ,
         \mem[43][5] , \mem[43][4] , \mem[43][3] , \mem[43][2] , \mem[43][1] ,
         \mem[43][0] , \mem[44][15] , \mem[44][14] , \mem[44][13] ,
         \mem[44][12] , \mem[44][11] , \mem[44][10] , \mem[44][9] ,
         \mem[44][8] , \mem[44][7] , \mem[44][6] , \mem[44][5] , \mem[44][4] ,
         \mem[44][3] , \mem[44][2] , \mem[44][1] , \mem[44][0] , \mem[45][15] ,
         \mem[45][14] , \mem[45][13] , \mem[45][12] , \mem[45][11] ,
         \mem[45][10] , \mem[45][9] , \mem[45][8] , \mem[45][7] , \mem[45][6] ,
         \mem[45][5] , \mem[45][4] , \mem[45][3] , \mem[45][2] , \mem[45][1] ,
         \mem[45][0] , \mem[46][15] , \mem[46][14] , \mem[46][13] ,
         \mem[46][12] , \mem[46][11] , \mem[46][10] , \mem[46][9] ,
         \mem[46][8] , \mem[46][7] , \mem[46][6] , \mem[46][5] , \mem[46][4] ,
         \mem[46][3] , \mem[46][2] , \mem[46][1] , \mem[46][0] , \mem[47][15] ,
         \mem[47][14] , \mem[47][13] , \mem[47][12] , \mem[47][11] ,
         \mem[47][10] , \mem[47][9] , \mem[47][8] , \mem[47][7] , \mem[47][6] ,
         \mem[47][5] , \mem[47][4] , \mem[47][3] , \mem[47][2] , \mem[47][1] ,
         \mem[47][0] , \mem[48][15] , \mem[48][14] , \mem[48][13] ,
         \mem[48][12] , \mem[48][11] , \mem[48][10] , \mem[48][9] ,
         \mem[48][8] , \mem[48][7] , \mem[48][6] , \mem[48][5] , \mem[48][4] ,
         \mem[48][3] , \mem[48][2] , \mem[48][1] , \mem[48][0] , \mem[49][15] ,
         \mem[49][14] , \mem[49][13] , \mem[49][12] , \mem[49][11] ,
         \mem[49][10] , \mem[49][9] , \mem[49][8] , \mem[49][7] , \mem[49][6] ,
         \mem[49][5] , \mem[49][4] , \mem[49][3] , \mem[49][2] , \mem[49][1] ,
         \mem[49][0] , \mem[50][15] , \mem[50][14] , \mem[50][13] ,
         \mem[50][12] , \mem[50][11] , \mem[50][10] , \mem[50][9] ,
         \mem[50][8] , \mem[50][7] , \mem[50][6] , \mem[50][5] , \mem[50][4] ,
         \mem[50][3] , \mem[50][2] , \mem[50][1] , \mem[50][0] , \mem[51][15] ,
         \mem[51][14] , \mem[51][13] , \mem[51][12] , \mem[51][11] ,
         \mem[51][10] , \mem[51][9] , \mem[51][8] , \mem[51][7] , \mem[51][6] ,
         \mem[51][5] , \mem[51][4] , \mem[51][3] , \mem[51][2] , \mem[51][1] ,
         \mem[51][0] , \mem[52][15] , \mem[52][14] , \mem[52][13] ,
         \mem[52][12] , \mem[52][11] , \mem[52][10] , \mem[52][9] ,
         \mem[52][8] , \mem[52][7] , \mem[52][6] , \mem[52][5] , \mem[52][4] ,
         \mem[52][3] , \mem[52][2] , \mem[52][1] , \mem[52][0] , \mem[53][15] ,
         \mem[53][14] , \mem[53][13] , \mem[53][12] , \mem[53][11] ,
         \mem[53][10] , \mem[53][9] , \mem[53][8] , \mem[53][7] , \mem[53][6] ,
         \mem[53][5] , \mem[53][4] , \mem[53][3] , \mem[53][2] , \mem[53][1] ,
         \mem[53][0] , \mem[54][15] , \mem[54][14] , \mem[54][13] ,
         \mem[54][12] , \mem[54][11] , \mem[54][10] , \mem[54][9] ,
         \mem[54][8] , \mem[54][7] , \mem[54][6] , \mem[54][5] , \mem[54][4] ,
         \mem[54][3] , \mem[54][2] , \mem[54][1] , \mem[54][0] , \mem[55][15] ,
         \mem[55][14] , \mem[55][13] , \mem[55][12] , \mem[55][11] ,
         \mem[55][10] , \mem[55][9] , \mem[55][8] , \mem[55][7] , \mem[55][6] ,
         \mem[55][5] , \mem[55][4] , \mem[55][3] , \mem[55][2] , \mem[55][1] ,
         \mem[55][0] , \mem[56][15] , \mem[56][14] , \mem[56][13] ,
         \mem[56][12] , \mem[56][11] , \mem[56][10] , \mem[56][9] ,
         \mem[56][8] , \mem[56][7] , \mem[56][6] , \mem[56][5] , \mem[56][4] ,
         \mem[56][3] , \mem[56][2] , \mem[56][1] , \mem[56][0] , \mem[57][15] ,
         \mem[57][14] , \mem[57][13] , \mem[57][12] , \mem[57][11] ,
         \mem[57][10] , \mem[57][9] , \mem[57][8] , \mem[57][7] , \mem[57][6] ,
         \mem[57][5] , \mem[57][4] , \mem[57][3] , \mem[57][2] , \mem[57][1] ,
         \mem[57][0] , \mem[58][15] , \mem[58][14] , \mem[58][13] ,
         \mem[58][12] , \mem[58][11] , \mem[58][10] , \mem[58][9] ,
         \mem[58][8] , \mem[58][7] , \mem[58][6] , \mem[58][5] , \mem[58][4] ,
         \mem[58][3] , \mem[58][2] , \mem[58][1] , \mem[58][0] , \mem[59][15] ,
         \mem[59][14] , \mem[59][13] , \mem[59][12] , \mem[59][11] ,
         \mem[59][10] , \mem[59][9] , \mem[59][8] , \mem[59][7] , \mem[59][6] ,
         \mem[59][5] , \mem[59][4] , \mem[59][3] , \mem[59][2] , \mem[59][1] ,
         \mem[59][0] , \mem[60][15] , \mem[60][14] , \mem[60][13] ,
         \mem[60][12] , \mem[60][11] , \mem[60][10] , \mem[60][9] ,
         \mem[60][8] , \mem[60][7] , \mem[60][6] , \mem[60][5] , \mem[60][4] ,
         \mem[60][3] , \mem[60][2] , \mem[60][1] , \mem[60][0] , \mem[61][15] ,
         \mem[61][14] , \mem[61][13] , \mem[61][12] , \mem[61][11] ,
         \mem[61][10] , \mem[61][9] , \mem[61][8] , \mem[61][7] , \mem[61][6] ,
         \mem[61][5] , \mem[61][4] , \mem[61][3] , \mem[61][2] , \mem[61][1] ,
         \mem[61][0] , \mem[62][15] , \mem[62][14] , \mem[62][13] ,
         \mem[62][12] , \mem[62][11] , \mem[62][10] , \mem[62][9] ,
         \mem[62][8] , \mem[62][7] , \mem[62][6] , \mem[62][5] , \mem[62][4] ,
         \mem[62][3] , \mem[62][2] , \mem[62][1] , \mem[62][0] , \mem[63][15] ,
         \mem[63][14] , \mem[63][13] , \mem[63][12] , \mem[63][11] ,
         \mem[63][10] , \mem[63][9] , \mem[63][8] , \mem[63][7] , \mem[63][6] ,
         \mem[63][5] , \mem[63][4] , \mem[63][3] , \mem[63][2] , \mem[63][1] ,
         \mem[63][0] , \mem[64][15] , \mem[64][14] , \mem[64][13] ,
         \mem[64][12] , \mem[64][11] , \mem[64][10] , \mem[64][9] ,
         \mem[64][8] , \mem[64][7] , \mem[64][6] , \mem[64][5] , \mem[64][4] ,
         \mem[64][3] , \mem[64][2] , \mem[64][1] , \mem[64][0] , \mem[65][15] ,
         \mem[65][14] , \mem[65][13] , \mem[65][12] , \mem[65][11] ,
         \mem[65][10] , \mem[65][9] , \mem[65][8] , \mem[65][7] , \mem[65][6] ,
         \mem[65][5] , \mem[65][4] , \mem[65][3] , \mem[65][2] , \mem[65][1] ,
         \mem[65][0] , \mem[66][15] , \mem[66][14] , \mem[66][13] ,
         \mem[66][12] , \mem[66][11] , \mem[66][10] , \mem[66][9] ,
         \mem[66][8] , \mem[66][7] , \mem[66][6] , \mem[66][5] , \mem[66][4] ,
         \mem[66][3] , \mem[66][2] , \mem[66][1] , \mem[66][0] , \mem[67][15] ,
         \mem[67][14] , \mem[67][13] , \mem[67][12] , \mem[67][11] ,
         \mem[67][10] , \mem[67][9] , \mem[67][8] , \mem[67][7] , \mem[67][6] ,
         \mem[67][5] , \mem[67][4] , \mem[67][3] , \mem[67][2] , \mem[67][1] ,
         \mem[67][0] , \mem[68][15] , \mem[68][14] , \mem[68][13] ,
         \mem[68][12] , \mem[68][11] , \mem[68][10] , \mem[68][9] ,
         \mem[68][8] , \mem[68][7] , \mem[68][6] , \mem[68][5] , \mem[68][4] ,
         \mem[68][3] , \mem[68][2] , \mem[68][1] , \mem[68][0] , \mem[69][15] ,
         \mem[69][14] , \mem[69][13] , \mem[69][12] , \mem[69][11] ,
         \mem[69][10] , \mem[69][9] , \mem[69][8] , \mem[69][7] , \mem[69][6] ,
         \mem[69][5] , \mem[69][4] , \mem[69][3] , \mem[69][2] , \mem[69][1] ,
         \mem[69][0] , \mem[70][15] , \mem[70][14] , \mem[70][13] ,
         \mem[70][12] , \mem[70][11] , \mem[70][10] , \mem[70][9] ,
         \mem[70][8] , \mem[70][7] , \mem[70][6] , \mem[70][5] , \mem[70][4] ,
         \mem[70][3] , \mem[70][2] , \mem[70][1] , \mem[70][0] , \mem[71][15] ,
         \mem[71][14] , \mem[71][13] , \mem[71][12] , \mem[71][11] ,
         \mem[71][10] , \mem[71][9] , \mem[71][8] , \mem[71][7] , \mem[71][6] ,
         \mem[71][5] , \mem[71][4] , \mem[71][3] , \mem[71][2] , \mem[71][1] ,
         \mem[71][0] , \mem[72][15] , \mem[72][14] , \mem[72][13] ,
         \mem[72][12] , \mem[72][11] , \mem[72][10] , \mem[72][9] ,
         \mem[72][8] , \mem[72][7] , \mem[72][6] , \mem[72][5] , \mem[72][4] ,
         \mem[72][3] , \mem[72][2] , \mem[72][1] , \mem[72][0] , \mem[73][15] ,
         \mem[73][14] , \mem[73][13] , \mem[73][12] , \mem[73][11] ,
         \mem[73][10] , \mem[73][9] , \mem[73][8] , \mem[73][7] , \mem[73][6] ,
         \mem[73][5] , \mem[73][4] , \mem[73][3] , \mem[73][2] , \mem[73][1] ,
         \mem[73][0] , \mem[74][15] , \mem[74][14] , \mem[74][13] ,
         \mem[74][12] , \mem[74][11] , \mem[74][10] , \mem[74][9] ,
         \mem[74][8] , \mem[74][7] , \mem[74][6] , \mem[74][5] , \mem[74][4] ,
         \mem[74][3] , \mem[74][2] , \mem[74][1] , \mem[74][0] , \mem[75][15] ,
         \mem[75][14] , \mem[75][13] , \mem[75][12] , \mem[75][11] ,
         \mem[75][10] , \mem[75][9] , \mem[75][8] , \mem[75][7] , \mem[75][6] ,
         \mem[75][5] , \mem[75][4] , \mem[75][3] , \mem[75][2] , \mem[75][1] ,
         \mem[75][0] , \mem[76][15] , \mem[76][14] , \mem[76][13] ,
         \mem[76][12] , \mem[76][11] , \mem[76][10] , \mem[76][9] ,
         \mem[76][8] , \mem[76][7] , \mem[76][6] , \mem[76][5] , \mem[76][4] ,
         \mem[76][3] , \mem[76][2] , \mem[76][1] , \mem[76][0] , \mem[77][15] ,
         \mem[77][14] , \mem[77][13] , \mem[77][12] , \mem[77][11] ,
         \mem[77][10] , \mem[77][9] , \mem[77][8] , \mem[77][7] , \mem[77][6] ,
         \mem[77][5] , \mem[77][4] , \mem[77][3] , \mem[77][2] , \mem[77][1] ,
         \mem[77][0] , \mem[78][15] , \mem[78][14] , \mem[78][13] ,
         \mem[78][12] , \mem[78][11] , \mem[78][10] , \mem[78][9] ,
         \mem[78][8] , \mem[78][7] , \mem[78][6] , \mem[78][5] , \mem[78][4] ,
         \mem[78][3] , \mem[78][2] , \mem[78][1] , \mem[78][0] , \mem[79][15] ,
         \mem[79][14] , \mem[79][13] , \mem[79][12] , \mem[79][11] ,
         \mem[79][10] , \mem[79][9] , \mem[79][8] , \mem[79][7] , \mem[79][6] ,
         \mem[79][5] , \mem[79][4] , \mem[79][3] , \mem[79][2] , \mem[79][1] ,
         \mem[79][0] , \mem[80][15] , \mem[80][14] , \mem[80][13] ,
         \mem[80][12] , \mem[80][11] , \mem[80][10] , \mem[80][9] ,
         \mem[80][8] , \mem[80][7] , \mem[80][6] , \mem[80][5] , \mem[80][4] ,
         \mem[80][3] , \mem[80][2] , \mem[80][1] , \mem[80][0] , \mem[81][15] ,
         \mem[81][14] , \mem[81][13] , \mem[81][12] , \mem[81][11] ,
         \mem[81][10] , \mem[81][9] , \mem[81][8] , \mem[81][7] , \mem[81][6] ,
         \mem[81][5] , \mem[81][4] , \mem[81][3] , \mem[81][2] , \mem[81][1] ,
         \mem[81][0] , \mem[82][15] , \mem[82][14] , \mem[82][13] ,
         \mem[82][12] , \mem[82][11] , \mem[82][10] , \mem[82][9] ,
         \mem[82][8] , \mem[82][7] , \mem[82][6] , \mem[82][5] , \mem[82][4] ,
         \mem[82][3] , \mem[82][2] , \mem[82][1] , \mem[82][0] , \mem[83][15] ,
         \mem[83][14] , \mem[83][13] , \mem[83][12] , \mem[83][11] ,
         \mem[83][10] , \mem[83][9] , \mem[83][8] , \mem[83][7] , \mem[83][6] ,
         \mem[83][5] , \mem[83][4] , \mem[83][3] , \mem[83][2] , \mem[83][1] ,
         \mem[83][0] , \mem[84][15] , \mem[84][14] , \mem[84][13] ,
         \mem[84][12] , \mem[84][11] , \mem[84][10] , \mem[84][9] ,
         \mem[84][8] , \mem[84][7] , \mem[84][6] , \mem[84][5] , \mem[84][4] ,
         \mem[84][3] , \mem[84][2] , \mem[84][1] , \mem[84][0] , \mem[85][15] ,
         \mem[85][14] , \mem[85][13] , \mem[85][12] , \mem[85][11] ,
         \mem[85][10] , \mem[85][9] , \mem[85][8] , \mem[85][7] , \mem[85][6] ,
         \mem[85][5] , \mem[85][4] , \mem[85][3] , \mem[85][2] , \mem[85][1] ,
         \mem[85][0] , \mem[86][15] , \mem[86][14] , \mem[86][13] ,
         \mem[86][12] , \mem[86][11] , \mem[86][10] , \mem[86][9] ,
         \mem[86][8] , \mem[86][7] , \mem[86][6] , \mem[86][5] , \mem[86][4] ,
         \mem[86][3] , \mem[86][2] , \mem[86][1] , \mem[86][0] , \mem[87][15] ,
         \mem[87][14] , \mem[87][13] , \mem[87][12] , \mem[87][11] ,
         \mem[87][10] , \mem[87][9] , \mem[87][8] , \mem[87][7] , \mem[87][6] ,
         \mem[87][5] , \mem[87][4] , \mem[87][3] , \mem[87][2] , \mem[87][1] ,
         \mem[87][0] , \mem[88][15] , \mem[88][14] , \mem[88][13] ,
         \mem[88][12] , \mem[88][11] , \mem[88][10] , \mem[88][9] ,
         \mem[88][8] , \mem[88][7] , \mem[88][6] , \mem[88][5] , \mem[88][4] ,
         \mem[88][3] , \mem[88][2] , \mem[88][1] , \mem[88][0] , \mem[89][15] ,
         \mem[89][14] , \mem[89][13] , \mem[89][12] , \mem[89][11] ,
         \mem[89][10] , \mem[89][9] , \mem[89][8] , \mem[89][7] , \mem[89][6] ,
         \mem[89][5] , \mem[89][4] , \mem[89][3] , \mem[89][2] , \mem[89][1] ,
         \mem[89][0] , \mem[90][15] , \mem[90][14] , \mem[90][13] ,
         \mem[90][12] , \mem[90][11] , \mem[90][10] , \mem[90][9] ,
         \mem[90][8] , \mem[90][7] , \mem[90][6] , \mem[90][5] , \mem[90][4] ,
         \mem[90][3] , \mem[90][2] , \mem[90][1] , \mem[90][0] , \mem[91][15] ,
         \mem[91][14] , \mem[91][13] , \mem[91][12] , \mem[91][11] ,
         \mem[91][10] , \mem[91][9] , \mem[91][8] , \mem[91][7] , \mem[91][6] ,
         \mem[91][5] , \mem[91][4] , \mem[91][3] , \mem[91][2] , \mem[91][1] ,
         \mem[91][0] , \mem[92][15] , \mem[92][14] , \mem[92][13] ,
         \mem[92][12] , \mem[92][11] , \mem[92][10] , \mem[92][9] ,
         \mem[92][8] , \mem[92][7] , \mem[92][6] , \mem[92][5] , \mem[92][4] ,
         \mem[92][3] , \mem[92][2] , \mem[92][1] , \mem[92][0] , \mem[93][15] ,
         \mem[93][14] , \mem[93][13] , \mem[93][12] , \mem[93][11] ,
         \mem[93][10] , \mem[93][9] , \mem[93][8] , \mem[93][7] , \mem[93][6] ,
         \mem[93][5] , \mem[93][4] , \mem[93][3] , \mem[93][2] , \mem[93][1] ,
         \mem[93][0] , \mem[94][15] , \mem[94][14] , \mem[94][13] ,
         \mem[94][12] , \mem[94][11] , \mem[94][10] , \mem[94][9] ,
         \mem[94][8] , \mem[94][7] , \mem[94][6] , \mem[94][5] , \mem[94][4] ,
         \mem[94][3] , \mem[94][2] , \mem[94][1] , \mem[94][0] , \mem[95][15] ,
         \mem[95][14] , \mem[95][13] , \mem[95][12] , \mem[95][11] ,
         \mem[95][10] , \mem[95][9] , \mem[95][8] , \mem[95][7] , \mem[95][6] ,
         \mem[95][5] , \mem[95][4] , \mem[95][3] , \mem[95][2] , \mem[95][1] ,
         \mem[95][0] , \mem[96][15] , \mem[96][14] , \mem[96][13] ,
         \mem[96][12] , \mem[96][11] , \mem[96][10] , \mem[96][9] ,
         \mem[96][8] , \mem[96][7] , \mem[96][6] , \mem[96][5] , \mem[96][4] ,
         \mem[96][3] , \mem[96][2] , \mem[96][1] , \mem[96][0] , \mem[97][15] ,
         \mem[97][14] , \mem[97][13] , \mem[97][12] , \mem[97][11] ,
         \mem[97][10] , \mem[97][9] , \mem[97][8] , \mem[97][7] , \mem[97][6] ,
         \mem[97][5] , \mem[97][4] , \mem[97][3] , \mem[97][2] , \mem[97][1] ,
         \mem[97][0] , \mem[98][15] , \mem[98][14] , \mem[98][13] ,
         \mem[98][12] , \mem[98][11] , \mem[98][10] , \mem[98][9] ,
         \mem[98][8] , \mem[98][7] , \mem[98][6] , \mem[98][5] , \mem[98][4] ,
         \mem[98][3] , \mem[98][2] , \mem[98][1] , \mem[98][0] , \mem[99][15] ,
         \mem[99][14] , \mem[99][13] , \mem[99][12] , \mem[99][11] ,
         \mem[99][10] , \mem[99][9] , \mem[99][8] , \mem[99][7] , \mem[99][6] ,
         \mem[99][5] , \mem[99][4] , \mem[99][3] , \mem[99][2] , \mem[99][1] ,
         \mem[99][0] , \mem[100][15] , \mem[100][14] , \mem[100][13] ,
         \mem[100][12] , \mem[100][11] , \mem[100][10] , \mem[100][9] ,
         \mem[100][8] , \mem[100][7] , \mem[100][6] , \mem[100][5] ,
         \mem[100][4] , \mem[100][3] , \mem[100][2] , \mem[100][1] ,
         \mem[100][0] , \mem[101][15] , \mem[101][14] , \mem[101][13] ,
         \mem[101][12] , \mem[101][11] , \mem[101][10] , \mem[101][9] ,
         \mem[101][8] , \mem[101][7] , \mem[101][6] , \mem[101][5] ,
         \mem[101][4] , \mem[101][3] , \mem[101][2] , \mem[101][1] ,
         \mem[101][0] , \mem[102][15] , \mem[102][14] , \mem[102][13] ,
         \mem[102][12] , \mem[102][11] , \mem[102][10] , \mem[102][9] ,
         \mem[102][8] , \mem[102][7] , \mem[102][6] , \mem[102][5] ,
         \mem[102][4] , \mem[102][3] , \mem[102][2] , \mem[102][1] ,
         \mem[102][0] , \mem[103][15] , \mem[103][14] , \mem[103][13] ,
         \mem[103][12] , \mem[103][11] , \mem[103][10] , \mem[103][9] ,
         \mem[103][8] , \mem[103][7] , \mem[103][6] , \mem[103][5] ,
         \mem[103][4] , \mem[103][3] , \mem[103][2] , \mem[103][1] ,
         \mem[103][0] , \mem[104][15] , \mem[104][14] , \mem[104][13] ,
         \mem[104][12] , \mem[104][11] , \mem[104][10] , \mem[104][9] ,
         \mem[104][8] , \mem[104][7] , \mem[104][6] , \mem[104][5] ,
         \mem[104][4] , \mem[104][3] , \mem[104][2] , \mem[104][1] ,
         \mem[104][0] , \mem[105][15] , \mem[105][14] , \mem[105][13] ,
         \mem[105][12] , \mem[105][11] , \mem[105][10] , \mem[105][9] ,
         \mem[105][8] , \mem[105][7] , \mem[105][6] , \mem[105][5] ,
         \mem[105][4] , \mem[105][3] , \mem[105][2] , \mem[105][1] ,
         \mem[105][0] , \mem[106][15] , \mem[106][14] , \mem[106][13] ,
         \mem[106][12] , \mem[106][11] , \mem[106][10] , \mem[106][9] ,
         \mem[106][8] , \mem[106][7] , \mem[106][6] , \mem[106][5] ,
         \mem[106][4] , \mem[106][3] , \mem[106][2] , \mem[106][1] ,
         \mem[106][0] , \mem[107][15] , \mem[107][14] , \mem[107][13] ,
         \mem[107][12] , \mem[107][11] , \mem[107][10] , \mem[107][9] ,
         \mem[107][8] , \mem[107][7] , \mem[107][6] , \mem[107][5] ,
         \mem[107][4] , \mem[107][3] , \mem[107][2] , \mem[107][1] ,
         \mem[107][0] , \mem[108][15] , \mem[108][14] , \mem[108][13] ,
         \mem[108][12] , \mem[108][11] , \mem[108][10] , \mem[108][9] ,
         \mem[108][8] , \mem[108][7] , \mem[108][6] , \mem[108][5] ,
         \mem[108][4] , \mem[108][3] , \mem[108][2] , \mem[108][1] ,
         \mem[108][0] , \mem[109][15] , \mem[109][14] , \mem[109][13] ,
         \mem[109][12] , \mem[109][11] , \mem[109][10] , \mem[109][9] ,
         \mem[109][8] , \mem[109][7] , \mem[109][6] , \mem[109][5] ,
         \mem[109][4] , \mem[109][3] , \mem[109][2] , \mem[109][1] ,
         \mem[109][0] , \mem[110][15] , \mem[110][14] , \mem[110][13] ,
         \mem[110][12] , \mem[110][11] , \mem[110][10] , \mem[110][9] ,
         \mem[110][8] , \mem[110][7] , \mem[110][6] , \mem[110][5] ,
         \mem[110][4] , \mem[110][3] , \mem[110][2] , \mem[110][1] ,
         \mem[110][0] , \mem[111][15] , \mem[111][14] , \mem[111][13] ,
         \mem[111][12] , \mem[111][11] , \mem[111][10] , \mem[111][9] ,
         \mem[111][8] , \mem[111][7] , \mem[111][6] , \mem[111][5] ,
         \mem[111][4] , \mem[111][3] , \mem[111][2] , \mem[111][1] ,
         \mem[111][0] , \mem[112][15] , \mem[112][14] , \mem[112][13] ,
         \mem[112][12] , \mem[112][11] , \mem[112][10] , \mem[112][9] ,
         \mem[112][8] , \mem[112][7] , \mem[112][6] , \mem[112][5] ,
         \mem[112][4] , \mem[112][3] , \mem[112][2] , \mem[112][1] ,
         \mem[112][0] , \mem[113][15] , \mem[113][14] , \mem[113][13] ,
         \mem[113][12] , \mem[113][11] , \mem[113][10] , \mem[113][9] ,
         \mem[113][8] , \mem[113][7] , \mem[113][6] , \mem[113][5] ,
         \mem[113][4] , \mem[113][3] , \mem[113][2] , \mem[113][1] ,
         \mem[113][0] , \mem[114][15] , \mem[114][14] , \mem[114][13] ,
         \mem[114][12] , \mem[114][11] , \mem[114][10] , \mem[114][9] ,
         \mem[114][8] , \mem[114][7] , \mem[114][6] , \mem[114][5] ,
         \mem[114][4] , \mem[114][3] , \mem[114][2] , \mem[114][1] ,
         \mem[114][0] , \mem[115][15] , \mem[115][14] , \mem[115][13] ,
         \mem[115][12] , \mem[115][11] , \mem[115][10] , \mem[115][9] ,
         \mem[115][8] , \mem[115][7] , \mem[115][6] , \mem[115][5] ,
         \mem[115][4] , \mem[115][3] , \mem[115][2] , \mem[115][1] ,
         \mem[115][0] , \mem[116][15] , \mem[116][14] , \mem[116][13] ,
         \mem[116][12] , \mem[116][11] , \mem[116][10] , \mem[116][9] ,
         \mem[116][8] , \mem[116][7] , \mem[116][6] , \mem[116][5] ,
         \mem[116][4] , \mem[116][3] , \mem[116][2] , \mem[116][1] ,
         \mem[116][0] , \mem[117][15] , \mem[117][14] , \mem[117][13] ,
         \mem[117][12] , \mem[117][11] , \mem[117][10] , \mem[117][9] ,
         \mem[117][8] , \mem[117][7] , \mem[117][6] , \mem[117][5] ,
         \mem[117][4] , \mem[117][3] , \mem[117][2] , \mem[117][1] ,
         \mem[117][0] , \mem[118][15] , \mem[118][14] , \mem[118][13] ,
         \mem[118][12] , \mem[118][11] , \mem[118][10] , \mem[118][9] ,
         \mem[118][8] , \mem[118][7] , \mem[118][6] , \mem[118][5] ,
         \mem[118][4] , \mem[118][3] , \mem[118][2] , \mem[118][1] ,
         \mem[118][0] , \mem[119][15] , \mem[119][14] , \mem[119][13] ,
         \mem[119][12] , \mem[119][11] , \mem[119][10] , \mem[119][9] ,
         \mem[119][8] , \mem[119][7] , \mem[119][6] , \mem[119][5] ,
         \mem[119][4] , \mem[119][3] , \mem[119][2] , \mem[119][1] ,
         \mem[119][0] , \mem[120][15] , \mem[120][14] , \mem[120][13] ,
         \mem[120][12] , \mem[120][11] , \mem[120][10] , \mem[120][9] ,
         \mem[120][8] , \mem[120][7] , \mem[120][6] , \mem[120][5] ,
         \mem[120][4] , \mem[120][3] , \mem[120][2] , \mem[120][1] ,
         \mem[120][0] , \mem[121][15] , \mem[121][14] , \mem[121][13] ,
         \mem[121][12] , \mem[121][11] , \mem[121][10] , \mem[121][9] ,
         \mem[121][8] , \mem[121][7] , \mem[121][6] , \mem[121][5] ,
         \mem[121][4] , \mem[121][3] , \mem[121][2] , \mem[121][1] ,
         \mem[121][0] , \mem[122][15] , \mem[122][14] , \mem[122][13] ,
         \mem[122][12] , \mem[122][11] , \mem[122][10] , \mem[122][9] ,
         \mem[122][8] , \mem[122][7] , \mem[122][6] , \mem[122][5] ,
         \mem[122][4] , \mem[122][3] , \mem[122][2] , \mem[122][1] ,
         \mem[122][0] , \mem[123][15] , \mem[123][14] , \mem[123][13] ,
         \mem[123][12] , \mem[123][11] , \mem[123][10] , \mem[123][9] ,
         \mem[123][8] , \mem[123][7] , \mem[123][6] , \mem[123][5] ,
         \mem[123][4] , \mem[123][3] , \mem[123][2] , \mem[123][1] ,
         \mem[123][0] , \mem[124][15] , \mem[124][14] , \mem[124][13] ,
         \mem[124][12] , \mem[124][11] , \mem[124][10] , \mem[124][9] ,
         \mem[124][8] , \mem[124][7] , \mem[124][6] , \mem[124][5] ,
         \mem[124][4] , \mem[124][3] , \mem[124][2] , \mem[124][1] ,
         \mem[124][0] , \mem[125][15] , \mem[125][14] , \mem[125][13] ,
         \mem[125][12] , \mem[125][11] , \mem[125][10] , \mem[125][9] ,
         \mem[125][8] , \mem[125][7] , \mem[125][6] , \mem[125][5] ,
         \mem[125][4] , \mem[125][3] , \mem[125][2] , \mem[125][1] ,
         \mem[125][0] , \mem[126][15] , \mem[126][14] , \mem[126][13] ,
         \mem[126][12] , \mem[126][11] , \mem[126][10] , \mem[126][9] ,
         \mem[126][8] , \mem[126][7] , \mem[126][6] , \mem[126][5] ,
         \mem[126][4] , \mem[126][3] , \mem[126][2] , \mem[126][1] ,
         \mem[126][0] , \mem[127][15] , \mem[127][14] , \mem[127][13] ,
         \mem[127][12] , \mem[127][11] , \mem[127][10] , \mem[127][9] ,
         \mem[127][8] , \mem[127][7] , \mem[127][6] , \mem[127][5] ,
         \mem[127][4] , \mem[127][3] , \mem[127][2] , \mem[127][1] ,
         \mem[127][0] , \mem[128][15] , \mem[128][14] , \mem[128][13] ,
         \mem[128][12] , \mem[128][11] , \mem[128][10] , \mem[128][9] ,
         \mem[128][8] , \mem[128][7] , \mem[128][6] , \mem[128][5] ,
         \mem[128][4] , \mem[128][3] , \mem[128][2] , \mem[128][1] ,
         \mem[128][0] , \mem[129][15] , \mem[129][14] , \mem[129][13] ,
         \mem[129][12] , \mem[129][11] , \mem[129][10] , \mem[129][9] ,
         \mem[129][8] , \mem[129][7] , \mem[129][6] , \mem[129][5] ,
         \mem[129][4] , \mem[129][3] , \mem[129][2] , \mem[129][1] ,
         \mem[129][0] , \mem[130][15] , \mem[130][14] , \mem[130][13] ,
         \mem[130][12] , \mem[130][11] , \mem[130][10] , \mem[130][9] ,
         \mem[130][8] , \mem[130][7] , \mem[130][6] , \mem[130][5] ,
         \mem[130][4] , \mem[130][3] , \mem[130][2] , \mem[130][1] ,
         \mem[130][0] , \mem[131][15] , \mem[131][14] , \mem[131][13] ,
         \mem[131][12] , \mem[131][11] , \mem[131][10] , \mem[131][9] ,
         \mem[131][8] , \mem[131][7] , \mem[131][6] , \mem[131][5] ,
         \mem[131][4] , \mem[131][3] , \mem[131][2] , \mem[131][1] ,
         \mem[131][0] , \mem[132][15] , \mem[132][14] , \mem[132][13] ,
         \mem[132][12] , \mem[132][11] , \mem[132][10] , \mem[132][9] ,
         \mem[132][8] , \mem[132][7] , \mem[132][6] , \mem[132][5] ,
         \mem[132][4] , \mem[132][3] , \mem[132][2] , \mem[132][1] ,
         \mem[132][0] , \mem[133][15] , \mem[133][14] , \mem[133][13] ,
         \mem[133][12] , \mem[133][11] , \mem[133][10] , \mem[133][9] ,
         \mem[133][8] , \mem[133][7] , \mem[133][6] , \mem[133][5] ,
         \mem[133][4] , \mem[133][3] , \mem[133][2] , \mem[133][1] ,
         \mem[133][0] , \mem[134][15] , \mem[134][14] , \mem[134][13] ,
         \mem[134][12] , \mem[134][11] , \mem[134][10] , \mem[134][9] ,
         \mem[134][8] , \mem[134][7] , \mem[134][6] , \mem[134][5] ,
         \mem[134][4] , \mem[134][3] , \mem[134][2] , \mem[134][1] ,
         \mem[134][0] , \mem[135][15] , \mem[135][14] , \mem[135][13] ,
         \mem[135][12] , \mem[135][11] , \mem[135][10] , \mem[135][9] ,
         \mem[135][8] , \mem[135][7] , \mem[135][6] , \mem[135][5] ,
         \mem[135][4] , \mem[135][3] , \mem[135][2] , \mem[135][1] ,
         \mem[135][0] , \mem[136][15] , \mem[136][14] , \mem[136][13] ,
         \mem[136][12] , \mem[136][11] , \mem[136][10] , \mem[136][9] ,
         \mem[136][8] , \mem[136][7] , \mem[136][6] , \mem[136][5] ,
         \mem[136][4] , \mem[136][3] , \mem[136][2] , \mem[136][1] ,
         \mem[136][0] , \mem[137][15] , \mem[137][14] , \mem[137][13] ,
         \mem[137][12] , \mem[137][11] , \mem[137][10] , \mem[137][9] ,
         \mem[137][8] , \mem[137][7] , \mem[137][6] , \mem[137][5] ,
         \mem[137][4] , \mem[137][3] , \mem[137][2] , \mem[137][1] ,
         \mem[137][0] , \mem[138][15] , \mem[138][14] , \mem[138][13] ,
         \mem[138][12] , \mem[138][11] , \mem[138][10] , \mem[138][9] ,
         \mem[138][8] , \mem[138][7] , \mem[138][6] , \mem[138][5] ,
         \mem[138][4] , \mem[138][3] , \mem[138][2] , \mem[138][1] ,
         \mem[138][0] , \mem[139][15] , \mem[139][14] , \mem[139][13] ,
         \mem[139][12] , \mem[139][11] , \mem[139][10] , \mem[139][9] ,
         \mem[139][8] , \mem[139][7] , \mem[139][6] , \mem[139][5] ,
         \mem[139][4] , \mem[139][3] , \mem[139][2] , \mem[139][1] ,
         \mem[139][0] , \mem[140][15] , \mem[140][14] , \mem[140][13] ,
         \mem[140][12] , \mem[140][11] , \mem[140][10] , \mem[140][9] ,
         \mem[140][8] , \mem[140][7] , \mem[140][6] , \mem[140][5] ,
         \mem[140][4] , \mem[140][3] , \mem[140][2] , \mem[140][1] ,
         \mem[140][0] , \mem[141][15] , \mem[141][14] , \mem[141][13] ,
         \mem[141][12] , \mem[141][11] , \mem[141][10] , \mem[141][9] ,
         \mem[141][8] , \mem[141][7] , \mem[141][6] , \mem[141][5] ,
         \mem[141][4] , \mem[141][3] , \mem[141][2] , \mem[141][1] ,
         \mem[141][0] , \mem[142][15] , \mem[142][14] , \mem[142][13] ,
         \mem[142][12] , \mem[142][11] , \mem[142][10] , \mem[142][9] ,
         \mem[142][8] , \mem[142][7] , \mem[142][6] , \mem[142][5] ,
         \mem[142][4] , \mem[142][3] , \mem[142][2] , \mem[142][1] ,
         \mem[142][0] , \mem[143][15] , \mem[143][14] , \mem[143][13] ,
         \mem[143][12] , \mem[143][11] , \mem[143][10] , \mem[143][9] ,
         \mem[143][8] , \mem[143][7] , \mem[143][6] , \mem[143][5] ,
         \mem[143][4] , \mem[143][3] , \mem[143][2] , \mem[143][1] ,
         \mem[143][0] , \mem[144][15] , \mem[144][14] , \mem[144][13] ,
         \mem[144][12] , \mem[144][11] , \mem[144][10] , \mem[144][9] ,
         \mem[144][8] , \mem[144][7] , \mem[144][6] , \mem[144][5] ,
         \mem[144][4] , \mem[144][3] , \mem[144][2] , \mem[144][1] ,
         \mem[144][0] , \mem[145][15] , \mem[145][14] , \mem[145][13] ,
         \mem[145][12] , \mem[145][11] , \mem[145][10] , \mem[145][9] ,
         \mem[145][8] , \mem[145][7] , \mem[145][6] , \mem[145][5] ,
         \mem[145][4] , \mem[145][3] , \mem[145][2] , \mem[145][1] ,
         \mem[145][0] , \mem[146][15] , \mem[146][14] , \mem[146][13] ,
         \mem[146][12] , \mem[146][11] , \mem[146][10] , \mem[146][9] ,
         \mem[146][8] , \mem[146][7] , \mem[146][6] , \mem[146][5] ,
         \mem[146][4] , \mem[146][3] , \mem[146][2] , \mem[146][1] ,
         \mem[146][0] , \mem[147][15] , \mem[147][14] , \mem[147][13] ,
         \mem[147][12] , \mem[147][11] , \mem[147][10] , \mem[147][9] ,
         \mem[147][8] , \mem[147][7] , \mem[147][6] , \mem[147][5] ,
         \mem[147][4] , \mem[147][3] , \mem[147][2] , \mem[147][1] ,
         \mem[147][0] , \mem[148][15] , \mem[148][14] , \mem[148][13] ,
         \mem[148][12] , \mem[148][11] , \mem[148][10] , \mem[148][9] ,
         \mem[148][8] , \mem[148][7] , \mem[148][6] , \mem[148][5] ,
         \mem[148][4] , \mem[148][3] , \mem[148][2] , \mem[148][1] ,
         \mem[148][0] , \mem[149][15] , \mem[149][14] , \mem[149][13] ,
         \mem[149][12] , \mem[149][11] , \mem[149][10] , \mem[149][9] ,
         \mem[149][8] , \mem[149][7] , \mem[149][6] , \mem[149][5] ,
         \mem[149][4] , \mem[149][3] , \mem[149][2] , \mem[149][1] ,
         \mem[149][0] , \mem[150][15] , \mem[150][14] , \mem[150][13] ,
         \mem[150][12] , \mem[150][11] , \mem[150][10] , \mem[150][9] ,
         \mem[150][8] , \mem[150][7] , \mem[150][6] , \mem[150][5] ,
         \mem[150][4] , \mem[150][3] , \mem[150][2] , \mem[150][1] ,
         \mem[150][0] , \mem[151][15] , \mem[151][14] , \mem[151][13] ,
         \mem[151][12] , \mem[151][11] , \mem[151][10] , \mem[151][9] ,
         \mem[151][8] , \mem[151][7] , \mem[151][6] , \mem[151][5] ,
         \mem[151][4] , \mem[151][3] , \mem[151][2] , \mem[151][1] ,
         \mem[151][0] , \mem[152][15] , \mem[152][14] , \mem[152][13] ,
         \mem[152][12] , \mem[152][11] , \mem[152][10] , \mem[152][9] ,
         \mem[152][8] , \mem[152][7] , \mem[152][6] , \mem[152][5] ,
         \mem[152][4] , \mem[152][3] , \mem[152][2] , \mem[152][1] ,
         \mem[152][0] , \mem[153][15] , \mem[153][14] , \mem[153][13] ,
         \mem[153][12] , \mem[153][11] , \mem[153][10] , \mem[153][9] ,
         \mem[153][8] , \mem[153][7] , \mem[153][6] , \mem[153][5] ,
         \mem[153][4] , \mem[153][3] , \mem[153][2] , \mem[153][1] ,
         \mem[153][0] , \mem[154][15] , \mem[154][14] , \mem[154][13] ,
         \mem[154][12] , \mem[154][11] , \mem[154][10] , \mem[154][9] ,
         \mem[154][8] , \mem[154][7] , \mem[154][6] , \mem[154][5] ,
         \mem[154][4] , \mem[154][3] , \mem[154][2] , \mem[154][1] ,
         \mem[154][0] , \mem[155][15] , \mem[155][14] , \mem[155][13] ,
         \mem[155][12] , \mem[155][11] , \mem[155][10] , \mem[155][9] ,
         \mem[155][8] , \mem[155][7] , \mem[155][6] , \mem[155][5] ,
         \mem[155][4] , \mem[155][3] , \mem[155][2] , \mem[155][1] ,
         \mem[155][0] , \mem[156][15] , \mem[156][14] , \mem[156][13] ,
         \mem[156][12] , \mem[156][11] , \mem[156][10] , \mem[156][9] ,
         \mem[156][8] , \mem[156][7] , \mem[156][6] , \mem[156][5] ,
         \mem[156][4] , \mem[156][3] , \mem[156][2] , \mem[156][1] ,
         \mem[156][0] , \mem[157][15] , \mem[157][14] , \mem[157][13] ,
         \mem[157][12] , \mem[157][11] , \mem[157][10] , \mem[157][9] ,
         \mem[157][8] , \mem[157][7] , \mem[157][6] , \mem[157][5] ,
         \mem[157][4] , \mem[157][3] , \mem[157][2] , \mem[157][1] ,
         \mem[157][0] , \mem[158][15] , \mem[158][14] , \mem[158][13] ,
         \mem[158][12] , \mem[158][11] , \mem[158][10] , \mem[158][9] ,
         \mem[158][8] , \mem[158][7] , \mem[158][6] , \mem[158][5] ,
         \mem[158][4] , \mem[158][3] , \mem[158][2] , \mem[158][1] ,
         \mem[158][0] , \mem[159][15] , \mem[159][14] , \mem[159][13] ,
         \mem[159][12] , \mem[159][11] , \mem[159][10] , \mem[159][9] ,
         \mem[159][8] , \mem[159][7] , \mem[159][6] , \mem[159][5] ,
         \mem[159][4] , \mem[159][3] , \mem[159][2] , \mem[159][1] ,
         \mem[159][0] , \mem[160][15] , \mem[160][14] , \mem[160][13] ,
         \mem[160][12] , \mem[160][11] , \mem[160][10] , \mem[160][9] ,
         \mem[160][8] , \mem[160][7] , \mem[160][6] , \mem[160][5] ,
         \mem[160][4] , \mem[160][3] , \mem[160][2] , \mem[160][1] ,
         \mem[160][0] , \mem[161][15] , \mem[161][14] , \mem[161][13] ,
         \mem[161][12] , \mem[161][11] , \mem[161][10] , \mem[161][9] ,
         \mem[161][8] , \mem[161][7] , \mem[161][6] , \mem[161][5] ,
         \mem[161][4] , \mem[161][3] , \mem[161][2] , \mem[161][1] ,
         \mem[161][0] , \mem[162][15] , \mem[162][14] , \mem[162][13] ,
         \mem[162][12] , \mem[162][11] , \mem[162][10] , \mem[162][9] ,
         \mem[162][8] , \mem[162][7] , \mem[162][6] , \mem[162][5] ,
         \mem[162][4] , \mem[162][3] , \mem[162][2] , \mem[162][1] ,
         \mem[162][0] , \mem[163][15] , \mem[163][14] , \mem[163][13] ,
         \mem[163][12] , \mem[163][11] , \mem[163][10] , \mem[163][9] ,
         \mem[163][8] , \mem[163][7] , \mem[163][6] , \mem[163][5] ,
         \mem[163][4] , \mem[163][3] , \mem[163][2] , \mem[163][1] ,
         \mem[163][0] , \mem[164][15] , \mem[164][14] , \mem[164][13] ,
         \mem[164][12] , \mem[164][11] , \mem[164][10] , \mem[164][9] ,
         \mem[164][8] , \mem[164][7] , \mem[164][6] , \mem[164][5] ,
         \mem[164][4] , \mem[164][3] , \mem[164][2] , \mem[164][1] ,
         \mem[164][0] , \mem[165][15] , \mem[165][14] , \mem[165][13] ,
         \mem[165][12] , \mem[165][11] , \mem[165][10] , \mem[165][9] ,
         \mem[165][8] , \mem[165][7] , \mem[165][6] , \mem[165][5] ,
         \mem[165][4] , \mem[165][3] , \mem[165][2] , \mem[165][1] ,
         \mem[165][0] , \mem[166][15] , \mem[166][14] , \mem[166][13] ,
         \mem[166][12] , \mem[166][11] , \mem[166][10] , \mem[166][9] ,
         \mem[166][8] , \mem[166][7] , \mem[166][6] , \mem[166][5] ,
         \mem[166][4] , \mem[166][3] , \mem[166][2] , \mem[166][1] ,
         \mem[166][0] , \mem[167][15] , \mem[167][14] , \mem[167][13] ,
         \mem[167][12] , \mem[167][11] , \mem[167][10] , \mem[167][9] ,
         \mem[167][8] , \mem[167][7] , \mem[167][6] , \mem[167][5] ,
         \mem[167][4] , \mem[167][3] , \mem[167][2] , \mem[167][1] ,
         \mem[167][0] , \mem[168][15] , \mem[168][14] , \mem[168][13] ,
         \mem[168][12] , \mem[168][11] , \mem[168][10] , \mem[168][9] ,
         \mem[168][8] , \mem[168][7] , \mem[168][6] , \mem[168][5] ,
         \mem[168][4] , \mem[168][3] , \mem[168][2] , \mem[168][1] ,
         \mem[168][0] , \mem[169][15] , \mem[169][14] , \mem[169][13] ,
         \mem[169][12] , \mem[169][11] , \mem[169][10] , \mem[169][9] ,
         \mem[169][8] , \mem[169][7] , \mem[169][6] , \mem[169][5] ,
         \mem[169][4] , \mem[169][3] , \mem[169][2] , \mem[169][1] ,
         \mem[169][0] , \mem[170][15] , \mem[170][14] , \mem[170][13] ,
         \mem[170][12] , \mem[170][11] , \mem[170][10] , \mem[170][9] ,
         \mem[170][8] , \mem[170][7] , \mem[170][6] , \mem[170][5] ,
         \mem[170][4] , \mem[170][3] , \mem[170][2] , \mem[170][1] ,
         \mem[170][0] , \mem[171][15] , \mem[171][14] , \mem[171][13] ,
         \mem[171][12] , \mem[171][11] , \mem[171][10] , \mem[171][9] ,
         \mem[171][8] , \mem[171][7] , \mem[171][6] , \mem[171][5] ,
         \mem[171][4] , \mem[171][3] , \mem[171][2] , \mem[171][1] ,
         \mem[171][0] , \mem[172][15] , \mem[172][14] , \mem[172][13] ,
         \mem[172][12] , \mem[172][11] , \mem[172][10] , \mem[172][9] ,
         \mem[172][8] , \mem[172][7] , \mem[172][6] , \mem[172][5] ,
         \mem[172][4] , \mem[172][3] , \mem[172][2] , \mem[172][1] ,
         \mem[172][0] , \mem[173][15] , \mem[173][14] , \mem[173][13] ,
         \mem[173][12] , \mem[173][11] , \mem[173][10] , \mem[173][9] ,
         \mem[173][8] , \mem[173][7] , \mem[173][6] , \mem[173][5] ,
         \mem[173][4] , \mem[173][3] , \mem[173][2] , \mem[173][1] ,
         \mem[173][0] , \mem[174][15] , \mem[174][14] , \mem[174][13] ,
         \mem[174][12] , \mem[174][11] , \mem[174][10] , \mem[174][9] ,
         \mem[174][8] , \mem[174][7] , \mem[174][6] , \mem[174][5] ,
         \mem[174][4] , \mem[174][3] , \mem[174][2] , \mem[174][1] ,
         \mem[174][0] , \mem[175][15] , \mem[175][14] , \mem[175][13] ,
         \mem[175][12] , \mem[175][11] , \mem[175][10] , \mem[175][9] ,
         \mem[175][8] , \mem[175][7] , \mem[175][6] , \mem[175][5] ,
         \mem[175][4] , \mem[175][3] , \mem[175][2] , \mem[175][1] ,
         \mem[175][0] , \mem[176][15] , \mem[176][14] , \mem[176][13] ,
         \mem[176][12] , \mem[176][11] , \mem[176][10] , \mem[176][9] ,
         \mem[176][8] , \mem[176][7] , \mem[176][6] , \mem[176][5] ,
         \mem[176][4] , \mem[176][3] , \mem[176][2] , \mem[176][1] ,
         \mem[176][0] , \mem[177][15] , \mem[177][14] , \mem[177][13] ,
         \mem[177][12] , \mem[177][11] , \mem[177][10] , \mem[177][9] ,
         \mem[177][8] , \mem[177][7] , \mem[177][6] , \mem[177][5] ,
         \mem[177][4] , \mem[177][3] , \mem[177][2] , \mem[177][1] ,
         \mem[177][0] , \mem[178][15] , \mem[178][14] , \mem[178][13] ,
         \mem[178][12] , \mem[178][11] , \mem[178][10] , \mem[178][9] ,
         \mem[178][8] , \mem[178][7] , \mem[178][6] , \mem[178][5] ,
         \mem[178][4] , \mem[178][3] , \mem[178][2] , \mem[178][1] ,
         \mem[178][0] , \mem[179][15] , \mem[179][14] , \mem[179][13] ,
         \mem[179][12] , \mem[179][11] , \mem[179][10] , \mem[179][9] ,
         \mem[179][8] , \mem[179][7] , \mem[179][6] , \mem[179][5] ,
         \mem[179][4] , \mem[179][3] , \mem[179][2] , \mem[179][1] ,
         \mem[179][0] , \mem[180][15] , \mem[180][14] , \mem[180][13] ,
         \mem[180][12] , \mem[180][11] , \mem[180][10] , \mem[180][9] ,
         \mem[180][8] , \mem[180][7] , \mem[180][6] , \mem[180][5] ,
         \mem[180][4] , \mem[180][3] , \mem[180][2] , \mem[180][1] ,
         \mem[180][0] , \mem[181][15] , \mem[181][14] , \mem[181][13] ,
         \mem[181][12] , \mem[181][11] , \mem[181][10] , \mem[181][9] ,
         \mem[181][8] , \mem[181][7] , \mem[181][6] , \mem[181][5] ,
         \mem[181][4] , \mem[181][3] , \mem[181][2] , \mem[181][1] ,
         \mem[181][0] , \mem[182][15] , \mem[182][14] , \mem[182][13] ,
         \mem[182][12] , \mem[182][11] , \mem[182][10] , \mem[182][9] ,
         \mem[182][8] , \mem[182][7] , \mem[182][6] , \mem[182][5] ,
         \mem[182][4] , \mem[182][3] , \mem[182][2] , \mem[182][1] ,
         \mem[182][0] , \mem[183][15] , \mem[183][14] , \mem[183][13] ,
         \mem[183][12] , \mem[183][11] , \mem[183][10] , \mem[183][9] ,
         \mem[183][8] , \mem[183][7] , \mem[183][6] , \mem[183][5] ,
         \mem[183][4] , \mem[183][3] , \mem[183][2] , \mem[183][1] ,
         \mem[183][0] , \mem[184][15] , \mem[184][14] , \mem[184][13] ,
         \mem[184][12] , \mem[184][11] , \mem[184][10] , \mem[184][9] ,
         \mem[184][8] , \mem[184][7] , \mem[184][6] , \mem[184][5] ,
         \mem[184][4] , \mem[184][3] , \mem[184][2] , \mem[184][1] ,
         \mem[184][0] , \mem[185][15] , \mem[185][14] , \mem[185][13] ,
         \mem[185][12] , \mem[185][11] , \mem[185][10] , \mem[185][9] ,
         \mem[185][8] , \mem[185][7] , \mem[185][6] , \mem[185][5] ,
         \mem[185][4] , \mem[185][3] , \mem[185][2] , \mem[185][1] ,
         \mem[185][0] , \mem[186][15] , \mem[186][14] , \mem[186][13] ,
         \mem[186][12] , \mem[186][11] , \mem[186][10] , \mem[186][9] ,
         \mem[186][8] , \mem[186][7] , \mem[186][6] , \mem[186][5] ,
         \mem[186][4] , \mem[186][3] , \mem[186][2] , \mem[186][1] ,
         \mem[186][0] , \mem[187][15] , \mem[187][14] , \mem[187][13] ,
         \mem[187][12] , \mem[187][11] , \mem[187][10] , \mem[187][9] ,
         \mem[187][8] , \mem[187][7] , \mem[187][6] , \mem[187][5] ,
         \mem[187][4] , \mem[187][3] , \mem[187][2] , \mem[187][1] ,
         \mem[187][0] , \mem[188][15] , \mem[188][14] , \mem[188][13] ,
         \mem[188][12] , \mem[188][11] , \mem[188][10] , \mem[188][9] ,
         \mem[188][8] , \mem[188][7] , \mem[188][6] , \mem[188][5] ,
         \mem[188][4] , \mem[188][3] , \mem[188][2] , \mem[188][1] ,
         \mem[188][0] , \mem[189][15] , \mem[189][14] , \mem[189][13] ,
         \mem[189][12] , \mem[189][11] , \mem[189][10] , \mem[189][9] ,
         \mem[189][8] , \mem[189][7] , \mem[189][6] , \mem[189][5] ,
         \mem[189][4] , \mem[189][3] , \mem[189][2] , \mem[189][1] ,
         \mem[189][0] , \mem[190][15] , \mem[190][14] , \mem[190][13] ,
         \mem[190][12] , \mem[190][11] , \mem[190][10] , \mem[190][9] ,
         \mem[190][8] , \mem[190][7] , \mem[190][6] , \mem[190][5] ,
         \mem[190][4] , \mem[190][3] , \mem[190][2] , \mem[190][1] ,
         \mem[190][0] , \mem[191][15] , \mem[191][14] , \mem[191][13] ,
         \mem[191][12] , \mem[191][11] , \mem[191][10] , \mem[191][9] ,
         \mem[191][8] , \mem[191][7] , \mem[191][6] , \mem[191][5] ,
         \mem[191][4] , \mem[191][3] , \mem[191][2] , \mem[191][1] ,
         \mem[191][0] , \mem[192][15] , \mem[192][14] , \mem[192][13] ,
         \mem[192][12] , \mem[192][11] , \mem[192][10] , \mem[192][9] ,
         \mem[192][8] , \mem[192][7] , \mem[192][6] , \mem[192][5] ,
         \mem[192][4] , \mem[192][3] , \mem[192][2] , \mem[192][1] ,
         \mem[192][0] , \mem[193][15] , \mem[193][14] , \mem[193][13] ,
         \mem[193][12] , \mem[193][11] , \mem[193][10] , \mem[193][9] ,
         \mem[193][8] , \mem[193][7] , \mem[193][6] , \mem[193][5] ,
         \mem[193][4] , \mem[193][3] , \mem[193][2] , \mem[193][1] ,
         \mem[193][0] , \mem[194][15] , \mem[194][14] , \mem[194][13] ,
         \mem[194][12] , \mem[194][11] , \mem[194][10] , \mem[194][9] ,
         \mem[194][8] , \mem[194][7] , \mem[194][6] , \mem[194][5] ,
         \mem[194][4] , \mem[194][3] , \mem[194][2] , \mem[194][1] ,
         \mem[194][0] , \mem[195][15] , \mem[195][14] , \mem[195][13] ,
         \mem[195][12] , \mem[195][11] , \mem[195][10] , \mem[195][9] ,
         \mem[195][8] , \mem[195][7] , \mem[195][6] , \mem[195][5] ,
         \mem[195][4] , \mem[195][3] , \mem[195][2] , \mem[195][1] ,
         \mem[195][0] , \mem[196][15] , \mem[196][14] , \mem[196][13] ,
         \mem[196][12] , \mem[196][11] , \mem[196][10] , \mem[196][9] ,
         \mem[196][8] , \mem[196][7] , \mem[196][6] , \mem[196][5] ,
         \mem[196][4] , \mem[196][3] , \mem[196][2] , \mem[196][1] ,
         \mem[196][0] , \mem[197][15] , \mem[197][14] , \mem[197][13] ,
         \mem[197][12] , \mem[197][11] , \mem[197][10] , \mem[197][9] ,
         \mem[197][8] , \mem[197][7] , \mem[197][6] , \mem[197][5] ,
         \mem[197][4] , \mem[197][3] , \mem[197][2] , \mem[197][1] ,
         \mem[197][0] , \mem[198][15] , \mem[198][14] , \mem[198][13] ,
         \mem[198][12] , \mem[198][11] , \mem[198][10] , \mem[198][9] ,
         \mem[198][8] , \mem[198][7] , \mem[198][6] , \mem[198][5] ,
         \mem[198][4] , \mem[198][3] , \mem[198][2] , \mem[198][1] ,
         \mem[198][0] , \mem[199][15] , \mem[199][14] , \mem[199][13] ,
         \mem[199][12] , \mem[199][11] , \mem[199][10] , \mem[199][9] ,
         \mem[199][8] , \mem[199][7] , \mem[199][6] , \mem[199][5] ,
         \mem[199][4] , \mem[199][3] , \mem[199][2] , \mem[199][1] ,
         \mem[199][0] , \mem[200][15] , \mem[200][14] , \mem[200][13] ,
         \mem[200][12] , \mem[200][11] , \mem[200][10] , \mem[200][9] ,
         \mem[200][8] , \mem[200][7] , \mem[200][6] , \mem[200][5] ,
         \mem[200][4] , \mem[200][3] , \mem[200][2] , \mem[200][1] ,
         \mem[200][0] , \mem[201][15] , \mem[201][14] , \mem[201][13] ,
         \mem[201][12] , \mem[201][11] , \mem[201][10] , \mem[201][9] ,
         \mem[201][8] , \mem[201][7] , \mem[201][6] , \mem[201][5] ,
         \mem[201][4] , \mem[201][3] , \mem[201][2] , \mem[201][1] ,
         \mem[201][0] , \mem[202][15] , \mem[202][14] , \mem[202][13] ,
         \mem[202][12] , \mem[202][11] , \mem[202][10] , \mem[202][9] ,
         \mem[202][8] , \mem[202][7] , \mem[202][6] , \mem[202][5] ,
         \mem[202][4] , \mem[202][3] , \mem[202][2] , \mem[202][1] ,
         \mem[202][0] , \mem[203][15] , \mem[203][14] , \mem[203][13] ,
         \mem[203][12] , \mem[203][11] , \mem[203][10] , \mem[203][9] ,
         \mem[203][8] , \mem[203][7] , \mem[203][6] , \mem[203][5] ,
         \mem[203][4] , \mem[203][3] , \mem[203][2] , \mem[203][1] ,
         \mem[203][0] , \mem[204][15] , \mem[204][14] , \mem[204][13] ,
         \mem[204][12] , \mem[204][11] , \mem[204][10] , \mem[204][9] ,
         \mem[204][8] , \mem[204][7] , \mem[204][6] , \mem[204][5] ,
         \mem[204][4] , \mem[204][3] , \mem[204][2] , \mem[204][1] ,
         \mem[204][0] , \mem[205][15] , \mem[205][14] , \mem[205][13] ,
         \mem[205][12] , \mem[205][11] , \mem[205][10] , \mem[205][9] ,
         \mem[205][8] , \mem[205][7] , \mem[205][6] , \mem[205][5] ,
         \mem[205][4] , \mem[205][3] , \mem[205][2] , \mem[205][1] ,
         \mem[205][0] , \mem[206][15] , \mem[206][14] , \mem[206][13] ,
         \mem[206][12] , \mem[206][11] , \mem[206][10] , \mem[206][9] ,
         \mem[206][8] , \mem[206][7] , \mem[206][6] , \mem[206][5] ,
         \mem[206][4] , \mem[206][3] , \mem[206][2] , \mem[206][1] ,
         \mem[206][0] , \mem[207][15] , \mem[207][14] , \mem[207][13] ,
         \mem[207][12] , \mem[207][11] , \mem[207][10] , \mem[207][9] ,
         \mem[207][8] , \mem[207][7] , \mem[207][6] , \mem[207][5] ,
         \mem[207][4] , \mem[207][3] , \mem[207][2] , \mem[207][1] ,
         \mem[207][0] , \mem[208][15] , \mem[208][14] , \mem[208][13] ,
         \mem[208][12] , \mem[208][11] , \mem[208][10] , \mem[208][9] ,
         \mem[208][8] , \mem[208][7] , \mem[208][6] , \mem[208][5] ,
         \mem[208][4] , \mem[208][3] , \mem[208][2] , \mem[208][1] ,
         \mem[208][0] , \mem[209][15] , \mem[209][14] , \mem[209][13] ,
         \mem[209][12] , \mem[209][11] , \mem[209][10] , \mem[209][9] ,
         \mem[209][8] , \mem[209][7] , \mem[209][6] , \mem[209][5] ,
         \mem[209][4] , \mem[209][3] , \mem[209][2] , \mem[209][1] ,
         \mem[209][0] , \mem[210][15] , \mem[210][14] , \mem[210][13] ,
         \mem[210][12] , \mem[210][11] , \mem[210][10] , \mem[210][9] ,
         \mem[210][8] , \mem[210][7] , \mem[210][6] , \mem[210][5] ,
         \mem[210][4] , \mem[210][3] , \mem[210][2] , \mem[210][1] ,
         \mem[210][0] , \mem[211][15] , \mem[211][14] , \mem[211][13] ,
         \mem[211][12] , \mem[211][11] , \mem[211][10] , \mem[211][9] ,
         \mem[211][8] , \mem[211][7] , \mem[211][6] , \mem[211][5] ,
         \mem[211][4] , \mem[211][3] , \mem[211][2] , \mem[211][1] ,
         \mem[211][0] , \mem[212][15] , \mem[212][14] , \mem[212][13] ,
         \mem[212][12] , \mem[212][11] , \mem[212][10] , \mem[212][9] ,
         \mem[212][8] , \mem[212][7] , \mem[212][6] , \mem[212][5] ,
         \mem[212][4] , \mem[212][3] , \mem[212][2] , \mem[212][1] ,
         \mem[212][0] , \mem[213][15] , \mem[213][14] , \mem[213][13] ,
         \mem[213][12] , \mem[213][11] , \mem[213][10] , \mem[213][9] ,
         \mem[213][8] , \mem[213][7] , \mem[213][6] , \mem[213][5] ,
         \mem[213][4] , \mem[213][3] , \mem[213][2] , \mem[213][1] ,
         \mem[213][0] , \mem[214][15] , \mem[214][14] , \mem[214][13] ,
         \mem[214][12] , \mem[214][11] , \mem[214][10] , \mem[214][9] ,
         \mem[214][8] , \mem[214][7] , \mem[214][6] , \mem[214][5] ,
         \mem[214][4] , \mem[214][3] , \mem[214][2] , \mem[214][1] ,
         \mem[214][0] , \mem[215][15] , \mem[215][14] , \mem[215][13] ,
         \mem[215][12] , \mem[215][11] , \mem[215][10] , \mem[215][9] ,
         \mem[215][8] , \mem[215][7] , \mem[215][6] , \mem[215][5] ,
         \mem[215][4] , \mem[215][3] , \mem[215][2] , \mem[215][1] ,
         \mem[215][0] , \mem[216][15] , \mem[216][14] , \mem[216][13] ,
         \mem[216][12] , \mem[216][11] , \mem[216][10] , \mem[216][9] ,
         \mem[216][8] , \mem[216][7] , \mem[216][6] , \mem[216][5] ,
         \mem[216][4] , \mem[216][3] , \mem[216][2] , \mem[216][1] ,
         \mem[216][0] , \mem[217][15] , \mem[217][14] , \mem[217][13] ,
         \mem[217][12] , \mem[217][11] , \mem[217][10] , \mem[217][9] ,
         \mem[217][8] , \mem[217][7] , \mem[217][6] , \mem[217][5] ,
         \mem[217][4] , \mem[217][3] , \mem[217][2] , \mem[217][1] ,
         \mem[217][0] , \mem[218][15] , \mem[218][14] , \mem[218][13] ,
         \mem[218][12] , \mem[218][11] , \mem[218][10] , \mem[218][9] ,
         \mem[218][8] , \mem[218][7] , \mem[218][6] , \mem[218][5] ,
         \mem[218][4] , \mem[218][3] , \mem[218][2] , \mem[218][1] ,
         \mem[218][0] , \mem[219][15] , \mem[219][14] , \mem[219][13] ,
         \mem[219][12] , \mem[219][11] , \mem[219][10] , \mem[219][9] ,
         \mem[219][8] , \mem[219][7] , \mem[219][6] , \mem[219][5] ,
         \mem[219][4] , \mem[219][3] , \mem[219][2] , \mem[219][1] ,
         \mem[219][0] , \mem[220][15] , \mem[220][14] , \mem[220][13] ,
         \mem[220][12] , \mem[220][11] , \mem[220][10] , \mem[220][9] ,
         \mem[220][8] , \mem[220][7] , \mem[220][6] , \mem[220][5] ,
         \mem[220][4] , \mem[220][3] , \mem[220][2] , \mem[220][1] ,
         \mem[220][0] , \mem[221][15] , \mem[221][14] , \mem[221][13] ,
         \mem[221][12] , \mem[221][11] , \mem[221][10] , \mem[221][9] ,
         \mem[221][8] , \mem[221][7] , \mem[221][6] , \mem[221][5] ,
         \mem[221][4] , \mem[221][3] , \mem[221][2] , \mem[221][1] ,
         \mem[221][0] , \mem[222][15] , \mem[222][14] , \mem[222][13] ,
         \mem[222][12] , \mem[222][11] , \mem[222][10] , \mem[222][9] ,
         \mem[222][8] , \mem[222][7] , \mem[222][6] , \mem[222][5] ,
         \mem[222][4] , \mem[222][3] , \mem[222][2] , \mem[222][1] ,
         \mem[222][0] , \mem[223][15] , \mem[223][14] , \mem[223][13] ,
         \mem[223][12] , \mem[223][11] , \mem[223][10] , \mem[223][9] ,
         \mem[223][8] , \mem[223][7] , \mem[223][6] , \mem[223][5] ,
         \mem[223][4] , \mem[223][3] , \mem[223][2] , \mem[223][1] ,
         \mem[223][0] , \mem[224][15] , \mem[224][14] , \mem[224][13] ,
         \mem[224][12] , \mem[224][11] , \mem[224][10] , \mem[224][9] ,
         \mem[224][8] , \mem[224][7] , \mem[224][6] , \mem[224][5] ,
         \mem[224][4] , \mem[224][3] , \mem[224][2] , \mem[224][1] ,
         \mem[224][0] , \mem[225][15] , \mem[225][14] , \mem[225][13] ,
         \mem[225][12] , \mem[225][11] , \mem[225][10] , \mem[225][9] ,
         \mem[225][8] , \mem[225][7] , \mem[225][6] , \mem[225][5] ,
         \mem[225][4] , \mem[225][3] , \mem[225][2] , \mem[225][1] ,
         \mem[225][0] , \mem[226][15] , \mem[226][14] , \mem[226][13] ,
         \mem[226][12] , \mem[226][11] , \mem[226][10] , \mem[226][9] ,
         \mem[226][8] , \mem[226][7] , \mem[226][6] , \mem[226][5] ,
         \mem[226][4] , \mem[226][3] , \mem[226][2] , \mem[226][1] ,
         \mem[226][0] , \mem[227][15] , \mem[227][14] , \mem[227][13] ,
         \mem[227][12] , \mem[227][11] , \mem[227][10] , \mem[227][9] ,
         \mem[227][8] , \mem[227][7] , \mem[227][6] , \mem[227][5] ,
         \mem[227][4] , \mem[227][3] , \mem[227][2] , \mem[227][1] ,
         \mem[227][0] , \mem[228][15] , \mem[228][14] , \mem[228][13] ,
         \mem[228][12] , \mem[228][11] , \mem[228][10] , \mem[228][9] ,
         \mem[228][8] , \mem[228][7] , \mem[228][6] , \mem[228][5] ,
         \mem[228][4] , \mem[228][3] , \mem[228][2] , \mem[228][1] ,
         \mem[228][0] , \mem[229][15] , \mem[229][14] , \mem[229][13] ,
         \mem[229][12] , \mem[229][11] , \mem[229][10] , \mem[229][9] ,
         \mem[229][8] , \mem[229][7] , \mem[229][6] , \mem[229][5] ,
         \mem[229][4] , \mem[229][3] , \mem[229][2] , \mem[229][1] ,
         \mem[229][0] , \mem[230][15] , \mem[230][14] , \mem[230][13] ,
         \mem[230][12] , \mem[230][11] , \mem[230][10] , \mem[230][9] ,
         \mem[230][8] , \mem[230][7] , \mem[230][6] , \mem[230][5] ,
         \mem[230][4] , \mem[230][3] , \mem[230][2] , \mem[230][1] ,
         \mem[230][0] , \mem[231][15] , \mem[231][14] , \mem[231][13] ,
         \mem[231][12] , \mem[231][11] , \mem[231][10] , \mem[231][9] ,
         \mem[231][8] , \mem[231][7] , \mem[231][6] , \mem[231][5] ,
         \mem[231][4] , \mem[231][3] , \mem[231][2] , \mem[231][1] ,
         \mem[231][0] , \mem[232][15] , \mem[232][14] , \mem[232][13] ,
         \mem[232][12] , \mem[232][11] , \mem[232][10] , \mem[232][9] ,
         \mem[232][8] , \mem[232][7] , \mem[232][6] , \mem[232][5] ,
         \mem[232][4] , \mem[232][3] , \mem[232][2] , \mem[232][1] ,
         \mem[232][0] , \mem[233][15] , \mem[233][14] , \mem[233][13] ,
         \mem[233][12] , \mem[233][11] , \mem[233][10] , \mem[233][9] ,
         \mem[233][8] , \mem[233][7] , \mem[233][6] , \mem[233][5] ,
         \mem[233][4] , \mem[233][3] , \mem[233][2] , \mem[233][1] ,
         \mem[233][0] , \mem[234][15] , \mem[234][14] , \mem[234][13] ,
         \mem[234][12] , \mem[234][11] , \mem[234][10] , \mem[234][9] ,
         \mem[234][8] , \mem[234][7] , \mem[234][6] , \mem[234][5] ,
         \mem[234][4] , \mem[234][3] , \mem[234][2] , \mem[234][1] ,
         \mem[234][0] , \mem[235][15] , \mem[235][14] , \mem[235][13] ,
         \mem[235][12] , \mem[235][11] , \mem[235][10] , \mem[235][9] ,
         \mem[235][8] , \mem[235][7] , \mem[235][6] , \mem[235][5] ,
         \mem[235][4] , \mem[235][3] , \mem[235][2] , \mem[235][1] ,
         \mem[235][0] , \mem[236][15] , \mem[236][14] , \mem[236][13] ,
         \mem[236][12] , \mem[236][11] , \mem[236][10] , \mem[236][9] ,
         \mem[236][8] , \mem[236][7] , \mem[236][6] , \mem[236][5] ,
         \mem[236][4] , \mem[236][3] , \mem[236][2] , \mem[236][1] ,
         \mem[236][0] , \mem[237][15] , \mem[237][14] , \mem[237][13] ,
         \mem[237][12] , \mem[237][11] , \mem[237][10] , \mem[237][9] ,
         \mem[237][8] , \mem[237][7] , \mem[237][6] , \mem[237][5] ,
         \mem[237][4] , \mem[237][3] , \mem[237][2] , \mem[237][1] ,
         \mem[237][0] , \mem[238][15] , \mem[238][14] , \mem[238][13] ,
         \mem[238][12] , \mem[238][11] , \mem[238][10] , \mem[238][9] ,
         \mem[238][8] , \mem[238][7] , \mem[238][6] , \mem[238][5] ,
         \mem[238][4] , \mem[238][3] , \mem[238][2] , \mem[238][1] ,
         \mem[238][0] , \mem[239][15] , \mem[239][14] , \mem[239][13] ,
         \mem[239][12] , \mem[239][11] , \mem[239][10] , \mem[239][9] ,
         \mem[239][8] , \mem[239][7] , \mem[239][6] , \mem[239][5] ,
         \mem[239][4] , \mem[239][3] , \mem[239][2] , \mem[239][1] ,
         \mem[239][0] , \mem[240][15] , \mem[240][14] , \mem[240][13] ,
         \mem[240][12] , \mem[240][11] , \mem[240][10] , \mem[240][9] ,
         \mem[240][8] , \mem[240][7] , \mem[240][6] , \mem[240][5] ,
         \mem[240][4] , \mem[240][3] , \mem[240][2] , \mem[240][1] ,
         \mem[240][0] , \mem[241][15] , \mem[241][14] , \mem[241][13] ,
         \mem[241][12] , \mem[241][11] , \mem[241][10] , \mem[241][9] ,
         \mem[241][8] , \mem[241][7] , \mem[241][6] , \mem[241][5] ,
         \mem[241][4] , \mem[241][3] , \mem[241][2] , \mem[241][1] ,
         \mem[241][0] , \mem[242][15] , \mem[242][14] , \mem[242][13] ,
         \mem[242][12] , \mem[242][11] , \mem[242][10] , \mem[242][9] ,
         \mem[242][8] , \mem[242][7] , \mem[242][6] , \mem[242][5] ,
         \mem[242][4] , \mem[242][3] , \mem[242][2] , \mem[242][1] ,
         \mem[242][0] , \mem[243][15] , \mem[243][14] , \mem[243][13] ,
         \mem[243][12] , \mem[243][11] , \mem[243][10] , \mem[243][9] ,
         \mem[243][8] , \mem[243][7] , \mem[243][6] , \mem[243][5] ,
         \mem[243][4] , \mem[243][3] , \mem[243][2] , \mem[243][1] ,
         \mem[243][0] , \mem[244][15] , \mem[244][14] , \mem[244][13] ,
         \mem[244][12] , \mem[244][11] , \mem[244][10] , \mem[244][9] ,
         \mem[244][8] , \mem[244][7] , \mem[244][6] , \mem[244][5] ,
         \mem[244][4] , \mem[244][3] , \mem[244][2] , \mem[244][1] ,
         \mem[244][0] , \mem[245][15] , \mem[245][14] , \mem[245][13] ,
         \mem[245][12] , \mem[245][11] , \mem[245][10] , \mem[245][9] ,
         \mem[245][8] , \mem[245][7] , \mem[245][6] , \mem[245][5] ,
         \mem[245][4] , \mem[245][3] , \mem[245][2] , \mem[245][1] ,
         \mem[245][0] , \mem[246][15] , \mem[246][14] , \mem[246][13] ,
         \mem[246][12] , \mem[246][11] , \mem[246][10] , \mem[246][9] ,
         \mem[246][8] , \mem[246][7] , \mem[246][6] , \mem[246][5] ,
         \mem[246][4] , \mem[246][3] , \mem[246][2] , \mem[246][1] ,
         \mem[246][0] , \mem[247][15] , \mem[247][14] , \mem[247][13] ,
         \mem[247][12] , \mem[247][11] , \mem[247][10] , \mem[247][9] ,
         \mem[247][8] , \mem[247][7] , \mem[247][6] , \mem[247][5] ,
         \mem[247][4] , \mem[247][3] , \mem[247][2] , \mem[247][1] ,
         \mem[247][0] , \mem[248][15] , \mem[248][14] , \mem[248][13] ,
         \mem[248][12] , \mem[248][11] , \mem[248][10] , \mem[248][9] ,
         \mem[248][8] , \mem[248][7] , \mem[248][6] , \mem[248][5] ,
         \mem[248][4] , \mem[248][3] , \mem[248][2] , \mem[248][1] ,
         \mem[248][0] , \mem[249][15] , \mem[249][14] , \mem[249][13] ,
         \mem[249][12] , \mem[249][11] , \mem[249][10] , \mem[249][9] ,
         \mem[249][8] , \mem[249][7] , \mem[249][6] , \mem[249][5] ,
         \mem[249][4] , \mem[249][3] , \mem[249][2] , \mem[249][1] ,
         \mem[249][0] , \mem[250][15] , \mem[250][14] , \mem[250][13] ,
         \mem[250][12] , \mem[250][11] , \mem[250][10] , \mem[250][9] ,
         \mem[250][8] , \mem[250][7] , \mem[250][6] , \mem[250][5] ,
         \mem[250][4] , \mem[250][3] , \mem[250][2] , \mem[250][1] ,
         \mem[250][0] , \mem[251][15] , \mem[251][14] , \mem[251][13] ,
         \mem[251][12] , \mem[251][11] , \mem[251][10] , \mem[251][9] ,
         \mem[251][8] , \mem[251][7] , \mem[251][6] , \mem[251][5] ,
         \mem[251][4] , \mem[251][3] , \mem[251][2] , \mem[251][1] ,
         \mem[251][0] , \mem[252][15] , \mem[252][14] , \mem[252][13] ,
         \mem[252][12] , \mem[252][11] , \mem[252][10] , \mem[252][9] ,
         \mem[252][8] , \mem[252][7] , \mem[252][6] , \mem[252][5] ,
         \mem[252][4] , \mem[252][3] , \mem[252][2] , \mem[252][1] ,
         \mem[252][0] , \mem[253][15] , \mem[253][14] , \mem[253][13] ,
         \mem[253][12] , \mem[253][11] , \mem[253][10] , \mem[253][9] ,
         \mem[253][8] , \mem[253][7] , \mem[253][6] , \mem[253][5] ,
         \mem[253][4] , \mem[253][3] , \mem[253][2] , \mem[253][1] ,
         \mem[253][0] , \mem[254][15] , \mem[254][14] , \mem[254][13] ,
         \mem[254][12] , \mem[254][11] , \mem[254][10] , \mem[254][9] ,
         \mem[254][8] , \mem[254][7] , \mem[254][6] , \mem[254][5] ,
         \mem[254][4] , \mem[254][3] , \mem[254][2] , \mem[254][1] ,
         \mem[254][0] , \mem[255][15] , \mem[255][14] , \mem[255][13] ,
         \mem[255][12] , \mem[255][11] , \mem[255][10] , \mem[255][9] ,
         \mem[255][8] , \mem[255][7] , \mem[255][6] , \mem[255][5] ,
         \mem[255][4] , \mem[255][3] , \mem[255][2] , \mem[255][1] ,
         \mem[255][0] , n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576;

  DFQD1 \mem_reg[0][15]  ( .D(n4668), .CP(clk), .Q(\mem[0][15] ) );
  DFQD1 \mem_reg[0][14]  ( .D(n4667), .CP(clk), .Q(\mem[0][14] ) );
  DFQD1 \mem_reg[0][13]  ( .D(n4666), .CP(clk), .Q(\mem[0][13] ) );
  DFQD1 \mem_reg[0][12]  ( .D(n4665), .CP(clk), .Q(\mem[0][12] ) );
  DFQD1 \mem_reg[0][11]  ( .D(n4664), .CP(clk), .Q(\mem[0][11] ) );
  DFQD1 \mem_reg[0][10]  ( .D(n4663), .CP(clk), .Q(\mem[0][10] ) );
  DFQD1 \mem_reg[0][9]  ( .D(n4662), .CP(clk), .Q(\mem[0][9] ) );
  DFQD1 \mem_reg[0][8]  ( .D(n4661), .CP(clk), .Q(\mem[0][8] ) );
  DFQD1 \mem_reg[0][7]  ( .D(n4660), .CP(clk), .Q(\mem[0][7] ) );
  DFQD1 \mem_reg[0][6]  ( .D(n4659), .CP(clk), .Q(\mem[0][6] ) );
  DFQD1 \mem_reg[0][5]  ( .D(n4658), .CP(clk), .Q(\mem[0][5] ) );
  DFQD1 \mem_reg[0][4]  ( .D(n4657), .CP(clk), .Q(\mem[0][4] ) );
  DFQD1 \mem_reg[0][3]  ( .D(n4656), .CP(clk), .Q(\mem[0][3] ) );
  DFQD1 \mem_reg[0][2]  ( .D(n4655), .CP(clk), .Q(\mem[0][2] ) );
  DFQD1 \mem_reg[0][1]  ( .D(n4654), .CP(clk), .Q(\mem[0][1] ) );
  DFQD1 \mem_reg[0][0]  ( .D(n4653), .CP(clk), .Q(\mem[0][0] ) );
  DFQD1 \mem_reg[1][15]  ( .D(n4652), .CP(clk), .Q(\mem[1][15] ) );
  DFQD1 \mem_reg[1][14]  ( .D(n4651), .CP(clk), .Q(\mem[1][14] ) );
  DFQD1 \mem_reg[1][13]  ( .D(n4650), .CP(clk), .Q(\mem[1][13] ) );
  DFQD1 \mem_reg[1][12]  ( .D(n4649), .CP(clk), .Q(\mem[1][12] ) );
  DFQD1 \mem_reg[1][11]  ( .D(n4648), .CP(clk), .Q(\mem[1][11] ) );
  DFQD1 \mem_reg[1][10]  ( .D(n4647), .CP(clk), .Q(\mem[1][10] ) );
  DFQD1 \mem_reg[1][9]  ( .D(n4646), .CP(clk), .Q(\mem[1][9] ) );
  DFQD1 \mem_reg[1][8]  ( .D(n4645), .CP(clk), .Q(\mem[1][8] ) );
  DFQD1 \mem_reg[1][7]  ( .D(n4644), .CP(clk), .Q(\mem[1][7] ) );
  DFQD1 \mem_reg[1][6]  ( .D(n4643), .CP(clk), .Q(\mem[1][6] ) );
  DFQD1 \mem_reg[1][5]  ( .D(n4642), .CP(clk), .Q(\mem[1][5] ) );
  DFQD1 \mem_reg[1][4]  ( .D(n4641), .CP(clk), .Q(\mem[1][4] ) );
  DFQD1 \mem_reg[1][3]  ( .D(n4640), .CP(clk), .Q(\mem[1][3] ) );
  DFQD1 \mem_reg[1][2]  ( .D(n4639), .CP(clk), .Q(\mem[1][2] ) );
  DFQD1 \mem_reg[1][1]  ( .D(n4638), .CP(clk), .Q(\mem[1][1] ) );
  DFQD1 \mem_reg[1][0]  ( .D(n4637), .CP(clk), .Q(\mem[1][0] ) );
  DFQD1 \mem_reg[2][15]  ( .D(n4636), .CP(clk), .Q(\mem[2][15] ) );
  DFQD1 \mem_reg[2][14]  ( .D(n4635), .CP(clk), .Q(\mem[2][14] ) );
  DFQD1 \mem_reg[2][13]  ( .D(n4634), .CP(clk), .Q(\mem[2][13] ) );
  DFQD1 \mem_reg[2][12]  ( .D(n4633), .CP(clk), .Q(\mem[2][12] ) );
  DFQD1 \mem_reg[2][11]  ( .D(n4632), .CP(clk), .Q(\mem[2][11] ) );
  DFQD1 \mem_reg[2][10]  ( .D(n4631), .CP(clk), .Q(\mem[2][10] ) );
  DFQD1 \mem_reg[2][9]  ( .D(n4630), .CP(clk), .Q(\mem[2][9] ) );
  DFQD1 \mem_reg[2][8]  ( .D(n4629), .CP(clk), .Q(\mem[2][8] ) );
  DFQD1 \mem_reg[2][7]  ( .D(n4628), .CP(clk), .Q(\mem[2][7] ) );
  DFQD1 \mem_reg[2][6]  ( .D(n4627), .CP(clk), .Q(\mem[2][6] ) );
  DFQD1 \mem_reg[2][5]  ( .D(n4626), .CP(clk), .Q(\mem[2][5] ) );
  DFQD1 \mem_reg[2][4]  ( .D(n4625), .CP(clk), .Q(\mem[2][4] ) );
  DFQD1 \mem_reg[2][3]  ( .D(n4624), .CP(clk), .Q(\mem[2][3] ) );
  DFQD1 \mem_reg[2][2]  ( .D(n4623), .CP(clk), .Q(\mem[2][2] ) );
  DFQD1 \mem_reg[2][1]  ( .D(n4622), .CP(clk), .Q(\mem[2][1] ) );
  DFQD1 \mem_reg[2][0]  ( .D(n4621), .CP(clk), .Q(\mem[2][0] ) );
  DFQD1 \mem_reg[3][15]  ( .D(n4620), .CP(clk), .Q(\mem[3][15] ) );
  DFQD1 \mem_reg[3][14]  ( .D(n4619), .CP(clk), .Q(\mem[3][14] ) );
  DFQD1 \mem_reg[3][13]  ( .D(n4618), .CP(clk), .Q(\mem[3][13] ) );
  DFQD1 \mem_reg[3][12]  ( .D(n4617), .CP(clk), .Q(\mem[3][12] ) );
  DFQD1 \mem_reg[3][11]  ( .D(n4616), .CP(clk), .Q(\mem[3][11] ) );
  DFQD1 \mem_reg[3][10]  ( .D(n4615), .CP(clk), .Q(\mem[3][10] ) );
  DFQD1 \mem_reg[3][9]  ( .D(n4614), .CP(clk), .Q(\mem[3][9] ) );
  DFQD1 \mem_reg[3][8]  ( .D(n4613), .CP(clk), .Q(\mem[3][8] ) );
  DFQD1 \mem_reg[3][7]  ( .D(n4612), .CP(clk), .Q(\mem[3][7] ) );
  DFQD1 \mem_reg[3][6]  ( .D(n4611), .CP(clk), .Q(\mem[3][6] ) );
  DFQD1 \mem_reg[3][5]  ( .D(n4610), .CP(clk), .Q(\mem[3][5] ) );
  DFQD1 \mem_reg[3][4]  ( .D(n4609), .CP(clk), .Q(\mem[3][4] ) );
  DFQD1 \mem_reg[3][3]  ( .D(n4608), .CP(clk), .Q(\mem[3][3] ) );
  DFQD1 \mem_reg[3][2]  ( .D(n4607), .CP(clk), .Q(\mem[3][2] ) );
  DFQD1 \mem_reg[3][1]  ( .D(n4606), .CP(clk), .Q(\mem[3][1] ) );
  DFQD1 \mem_reg[3][0]  ( .D(n4605), .CP(clk), .Q(\mem[3][0] ) );
  DFQD1 \mem_reg[4][15]  ( .D(n4604), .CP(clk), .Q(\mem[4][15] ) );
  DFQD1 \mem_reg[4][14]  ( .D(n4603), .CP(clk), .Q(\mem[4][14] ) );
  DFQD1 \mem_reg[4][13]  ( .D(n4602), .CP(clk), .Q(\mem[4][13] ) );
  DFQD1 \mem_reg[4][12]  ( .D(n4601), .CP(clk), .Q(\mem[4][12] ) );
  DFQD1 \mem_reg[4][11]  ( .D(n4600), .CP(clk), .Q(\mem[4][11] ) );
  DFQD1 \mem_reg[4][10]  ( .D(n4599), .CP(clk), .Q(\mem[4][10] ) );
  DFQD1 \mem_reg[4][9]  ( .D(n4598), .CP(clk), .Q(\mem[4][9] ) );
  DFQD1 \mem_reg[4][8]  ( .D(n4597), .CP(clk), .Q(\mem[4][8] ) );
  DFQD1 \mem_reg[4][7]  ( .D(n4596), .CP(clk), .Q(\mem[4][7] ) );
  DFQD1 \mem_reg[4][6]  ( .D(n4595), .CP(clk), .Q(\mem[4][6] ) );
  DFQD1 \mem_reg[4][5]  ( .D(n4594), .CP(clk), .Q(\mem[4][5] ) );
  DFQD1 \mem_reg[4][4]  ( .D(n4593), .CP(clk), .Q(\mem[4][4] ) );
  DFQD1 \mem_reg[4][3]  ( .D(n4592), .CP(clk), .Q(\mem[4][3] ) );
  DFQD1 \mem_reg[4][2]  ( .D(n4591), .CP(clk), .Q(\mem[4][2] ) );
  DFQD1 \mem_reg[4][1]  ( .D(n4590), .CP(clk), .Q(\mem[4][1] ) );
  DFQD1 \mem_reg[4][0]  ( .D(n4589), .CP(clk), .Q(\mem[4][0] ) );
  DFQD1 \mem_reg[5][15]  ( .D(n4588), .CP(clk), .Q(\mem[5][15] ) );
  DFQD1 \mem_reg[5][14]  ( .D(n4587), .CP(clk), .Q(\mem[5][14] ) );
  DFQD1 \mem_reg[5][13]  ( .D(n4586), .CP(clk), .Q(\mem[5][13] ) );
  DFQD1 \mem_reg[5][12]  ( .D(n4585), .CP(clk), .Q(\mem[5][12] ) );
  DFQD1 \mem_reg[5][11]  ( .D(n4584), .CP(clk), .Q(\mem[5][11] ) );
  DFQD1 \mem_reg[5][10]  ( .D(n4583), .CP(clk), .Q(\mem[5][10] ) );
  DFQD1 \mem_reg[5][9]  ( .D(n4582), .CP(clk), .Q(\mem[5][9] ) );
  DFQD1 \mem_reg[5][8]  ( .D(n4581), .CP(clk), .Q(\mem[5][8] ) );
  DFQD1 \mem_reg[5][7]  ( .D(n4580), .CP(clk), .Q(\mem[5][7] ) );
  DFQD1 \mem_reg[5][6]  ( .D(n4579), .CP(clk), .Q(\mem[5][6] ) );
  DFQD1 \mem_reg[5][5]  ( .D(n4578), .CP(clk), .Q(\mem[5][5] ) );
  DFQD1 \mem_reg[5][4]  ( .D(n4577), .CP(clk), .Q(\mem[5][4] ) );
  DFQD1 \mem_reg[5][3]  ( .D(n4576), .CP(clk), .Q(\mem[5][3] ) );
  DFQD1 \mem_reg[5][2]  ( .D(n4575), .CP(clk), .Q(\mem[5][2] ) );
  DFQD1 \mem_reg[5][1]  ( .D(n4574), .CP(clk), .Q(\mem[5][1] ) );
  DFQD1 \mem_reg[5][0]  ( .D(n4573), .CP(clk), .Q(\mem[5][0] ) );
  DFQD1 \mem_reg[6][15]  ( .D(n4572), .CP(clk), .Q(\mem[6][15] ) );
  DFQD1 \mem_reg[6][14]  ( .D(n4571), .CP(clk), .Q(\mem[6][14] ) );
  DFQD1 \mem_reg[6][13]  ( .D(n4570), .CP(clk), .Q(\mem[6][13] ) );
  DFQD1 \mem_reg[6][12]  ( .D(n4569), .CP(clk), .Q(\mem[6][12] ) );
  DFQD1 \mem_reg[6][11]  ( .D(n4568), .CP(clk), .Q(\mem[6][11] ) );
  DFQD1 \mem_reg[6][10]  ( .D(n4567), .CP(clk), .Q(\mem[6][10] ) );
  DFQD1 \mem_reg[6][9]  ( .D(n4566), .CP(clk), .Q(\mem[6][9] ) );
  DFQD1 \mem_reg[6][8]  ( .D(n4565), .CP(clk), .Q(\mem[6][8] ) );
  DFQD1 \mem_reg[6][7]  ( .D(n4564), .CP(clk), .Q(\mem[6][7] ) );
  DFQD1 \mem_reg[6][6]  ( .D(n4563), .CP(clk), .Q(\mem[6][6] ) );
  DFQD1 \mem_reg[6][5]  ( .D(n4562), .CP(clk), .Q(\mem[6][5] ) );
  DFQD1 \mem_reg[6][4]  ( .D(n4561), .CP(clk), .Q(\mem[6][4] ) );
  DFQD1 \mem_reg[6][3]  ( .D(n4560), .CP(clk), .Q(\mem[6][3] ) );
  DFQD1 \mem_reg[6][2]  ( .D(n4559), .CP(clk), .Q(\mem[6][2] ) );
  DFQD1 \mem_reg[6][1]  ( .D(n4558), .CP(clk), .Q(\mem[6][1] ) );
  DFQD1 \mem_reg[6][0]  ( .D(n4557), .CP(clk), .Q(\mem[6][0] ) );
  DFQD1 \mem_reg[7][15]  ( .D(n4556), .CP(clk), .Q(\mem[7][15] ) );
  DFQD1 \mem_reg[7][14]  ( .D(n4555), .CP(clk), .Q(\mem[7][14] ) );
  DFQD1 \mem_reg[7][13]  ( .D(n4554), .CP(clk), .Q(\mem[7][13] ) );
  DFQD1 \mem_reg[7][12]  ( .D(n4553), .CP(clk), .Q(\mem[7][12] ) );
  DFQD1 \mem_reg[7][11]  ( .D(n4552), .CP(clk), .Q(\mem[7][11] ) );
  DFQD1 \mem_reg[7][10]  ( .D(n4551), .CP(clk), .Q(\mem[7][10] ) );
  DFQD1 \mem_reg[7][9]  ( .D(n4550), .CP(clk), .Q(\mem[7][9] ) );
  DFQD1 \mem_reg[7][8]  ( .D(n4549), .CP(clk), .Q(\mem[7][8] ) );
  DFQD1 \mem_reg[7][7]  ( .D(n4548), .CP(clk), .Q(\mem[7][7] ) );
  DFQD1 \mem_reg[7][6]  ( .D(n4547), .CP(clk), .Q(\mem[7][6] ) );
  DFQD1 \mem_reg[7][5]  ( .D(n4546), .CP(clk), .Q(\mem[7][5] ) );
  DFQD1 \mem_reg[7][4]  ( .D(n4545), .CP(clk), .Q(\mem[7][4] ) );
  DFQD1 \mem_reg[7][3]  ( .D(n4544), .CP(clk), .Q(\mem[7][3] ) );
  DFQD1 \mem_reg[7][2]  ( .D(n4543), .CP(clk), .Q(\mem[7][2] ) );
  DFQD1 \mem_reg[7][1]  ( .D(n4542), .CP(clk), .Q(\mem[7][1] ) );
  DFQD1 \mem_reg[7][0]  ( .D(n4541), .CP(clk), .Q(\mem[7][0] ) );
  DFQD1 \mem_reg[8][15]  ( .D(n4540), .CP(clk), .Q(\mem[8][15] ) );
  DFQD1 \mem_reg[8][14]  ( .D(n4539), .CP(clk), .Q(\mem[8][14] ) );
  DFQD1 \mem_reg[8][13]  ( .D(n4538), .CP(clk), .Q(\mem[8][13] ) );
  DFQD1 \mem_reg[8][12]  ( .D(n4537), .CP(clk), .Q(\mem[8][12] ) );
  DFQD1 \mem_reg[8][11]  ( .D(n4536), .CP(clk), .Q(\mem[8][11] ) );
  DFQD1 \mem_reg[8][10]  ( .D(n4535), .CP(clk), .Q(\mem[8][10] ) );
  DFQD1 \mem_reg[8][9]  ( .D(n4534), .CP(clk), .Q(\mem[8][9] ) );
  DFQD1 \mem_reg[8][8]  ( .D(n4533), .CP(clk), .Q(\mem[8][8] ) );
  DFQD1 \mem_reg[8][7]  ( .D(n4532), .CP(clk), .Q(\mem[8][7] ) );
  DFQD1 \mem_reg[8][6]  ( .D(n4531), .CP(clk), .Q(\mem[8][6] ) );
  DFQD1 \mem_reg[8][5]  ( .D(n4530), .CP(clk), .Q(\mem[8][5] ) );
  DFQD1 \mem_reg[8][4]  ( .D(n4529), .CP(clk), .Q(\mem[8][4] ) );
  DFQD1 \mem_reg[8][3]  ( .D(n4528), .CP(clk), .Q(\mem[8][3] ) );
  DFQD1 \mem_reg[8][2]  ( .D(n4527), .CP(clk), .Q(\mem[8][2] ) );
  DFQD1 \mem_reg[8][1]  ( .D(n4526), .CP(clk), .Q(\mem[8][1] ) );
  DFQD1 \mem_reg[8][0]  ( .D(n4525), .CP(clk), .Q(\mem[8][0] ) );
  DFQD1 \mem_reg[9][15]  ( .D(n4524), .CP(clk), .Q(\mem[9][15] ) );
  DFQD1 \mem_reg[9][14]  ( .D(n4523), .CP(clk), .Q(\mem[9][14] ) );
  DFQD1 \mem_reg[9][13]  ( .D(n4522), .CP(clk), .Q(\mem[9][13] ) );
  DFQD1 \mem_reg[9][12]  ( .D(n4521), .CP(clk), .Q(\mem[9][12] ) );
  DFQD1 \mem_reg[9][11]  ( .D(n4520), .CP(clk), .Q(\mem[9][11] ) );
  DFQD1 \mem_reg[9][10]  ( .D(n4519), .CP(clk), .Q(\mem[9][10] ) );
  DFQD1 \mem_reg[9][9]  ( .D(n4518), .CP(clk), .Q(\mem[9][9] ) );
  DFQD1 \mem_reg[9][8]  ( .D(n4517), .CP(clk), .Q(\mem[9][8] ) );
  DFQD1 \mem_reg[9][7]  ( .D(n4516), .CP(clk), .Q(\mem[9][7] ) );
  DFQD1 \mem_reg[9][6]  ( .D(n4515), .CP(clk), .Q(\mem[9][6] ) );
  DFQD1 \mem_reg[9][5]  ( .D(n4514), .CP(clk), .Q(\mem[9][5] ) );
  DFQD1 \mem_reg[9][4]  ( .D(n4513), .CP(clk), .Q(\mem[9][4] ) );
  DFQD1 \mem_reg[9][3]  ( .D(n4512), .CP(clk), .Q(\mem[9][3] ) );
  DFQD1 \mem_reg[9][2]  ( .D(n4511), .CP(clk), .Q(\mem[9][2] ) );
  DFQD1 \mem_reg[9][1]  ( .D(n4510), .CP(clk), .Q(\mem[9][1] ) );
  DFQD1 \mem_reg[9][0]  ( .D(n4509), .CP(clk), .Q(\mem[9][0] ) );
  DFQD1 \mem_reg[10][15]  ( .D(n4508), .CP(clk), .Q(\mem[10][15] ) );
  DFQD1 \mem_reg[10][14]  ( .D(n4507), .CP(clk), .Q(\mem[10][14] ) );
  DFQD1 \mem_reg[10][13]  ( .D(n4506), .CP(clk), .Q(\mem[10][13] ) );
  DFQD1 \mem_reg[10][12]  ( .D(n4505), .CP(clk), .Q(\mem[10][12] ) );
  DFQD1 \mem_reg[10][11]  ( .D(n4504), .CP(clk), .Q(\mem[10][11] ) );
  DFQD1 \mem_reg[10][10]  ( .D(n4503), .CP(clk), .Q(\mem[10][10] ) );
  DFQD1 \mem_reg[10][9]  ( .D(n4502), .CP(clk), .Q(\mem[10][9] ) );
  DFQD1 \mem_reg[10][8]  ( .D(n4501), .CP(clk), .Q(\mem[10][8] ) );
  DFQD1 \mem_reg[10][7]  ( .D(n4500), .CP(clk), .Q(\mem[10][7] ) );
  DFQD1 \mem_reg[10][6]  ( .D(n4499), .CP(clk), .Q(\mem[10][6] ) );
  DFQD1 \mem_reg[10][5]  ( .D(n4498), .CP(clk), .Q(\mem[10][5] ) );
  DFQD1 \mem_reg[10][4]  ( .D(n4497), .CP(clk), .Q(\mem[10][4] ) );
  DFQD1 \mem_reg[10][3]  ( .D(n4496), .CP(clk), .Q(\mem[10][3] ) );
  DFQD1 \mem_reg[10][2]  ( .D(n4495), .CP(clk), .Q(\mem[10][2] ) );
  DFQD1 \mem_reg[10][1]  ( .D(n4494), .CP(clk), .Q(\mem[10][1] ) );
  DFQD1 \mem_reg[10][0]  ( .D(n4493), .CP(clk), .Q(\mem[10][0] ) );
  DFQD1 \mem_reg[11][15]  ( .D(n4492), .CP(clk), .Q(\mem[11][15] ) );
  DFQD1 \mem_reg[11][14]  ( .D(n4491), .CP(clk), .Q(\mem[11][14] ) );
  DFQD1 \mem_reg[11][13]  ( .D(n4490), .CP(clk), .Q(\mem[11][13] ) );
  DFQD1 \mem_reg[11][12]  ( .D(n4489), .CP(clk), .Q(\mem[11][12] ) );
  DFQD1 \mem_reg[11][11]  ( .D(n4488), .CP(clk), .Q(\mem[11][11] ) );
  DFQD1 \mem_reg[11][10]  ( .D(n4487), .CP(clk), .Q(\mem[11][10] ) );
  DFQD1 \mem_reg[11][9]  ( .D(n4486), .CP(clk), .Q(\mem[11][9] ) );
  DFQD1 \mem_reg[11][8]  ( .D(n4485), .CP(clk), .Q(\mem[11][8] ) );
  DFQD1 \mem_reg[11][7]  ( .D(n4484), .CP(clk), .Q(\mem[11][7] ) );
  DFQD1 \mem_reg[11][6]  ( .D(n4483), .CP(clk), .Q(\mem[11][6] ) );
  DFQD1 \mem_reg[11][5]  ( .D(n4482), .CP(clk), .Q(\mem[11][5] ) );
  DFQD1 \mem_reg[11][4]  ( .D(n4481), .CP(clk), .Q(\mem[11][4] ) );
  DFQD1 \mem_reg[11][3]  ( .D(n4480), .CP(clk), .Q(\mem[11][3] ) );
  DFQD1 \mem_reg[11][2]  ( .D(n4479), .CP(clk), .Q(\mem[11][2] ) );
  DFQD1 \mem_reg[11][1]  ( .D(n4478), .CP(clk), .Q(\mem[11][1] ) );
  DFQD1 \mem_reg[11][0]  ( .D(n4477), .CP(clk), .Q(\mem[11][0] ) );
  DFQD1 \mem_reg[12][15]  ( .D(n4476), .CP(clk), .Q(\mem[12][15] ) );
  DFQD1 \mem_reg[12][14]  ( .D(n4475), .CP(clk), .Q(\mem[12][14] ) );
  DFQD1 \mem_reg[12][13]  ( .D(n4474), .CP(clk), .Q(\mem[12][13] ) );
  DFQD1 \mem_reg[12][12]  ( .D(n4473), .CP(clk), .Q(\mem[12][12] ) );
  DFQD1 \mem_reg[12][11]  ( .D(n4472), .CP(clk), .Q(\mem[12][11] ) );
  DFQD1 \mem_reg[12][10]  ( .D(n4471), .CP(clk), .Q(\mem[12][10] ) );
  DFQD1 \mem_reg[12][9]  ( .D(n4470), .CP(clk), .Q(\mem[12][9] ) );
  DFQD1 \mem_reg[12][8]  ( .D(n4469), .CP(clk), .Q(\mem[12][8] ) );
  DFQD1 \mem_reg[12][7]  ( .D(n4468), .CP(clk), .Q(\mem[12][7] ) );
  DFQD1 \mem_reg[12][6]  ( .D(n4467), .CP(clk), .Q(\mem[12][6] ) );
  DFQD1 \mem_reg[12][5]  ( .D(n4466), .CP(clk), .Q(\mem[12][5] ) );
  DFQD1 \mem_reg[12][4]  ( .D(n4465), .CP(clk), .Q(\mem[12][4] ) );
  DFQD1 \mem_reg[12][3]  ( .D(n4464), .CP(clk), .Q(\mem[12][3] ) );
  DFQD1 \mem_reg[12][2]  ( .D(n4463), .CP(clk), .Q(\mem[12][2] ) );
  DFQD1 \mem_reg[12][1]  ( .D(n4462), .CP(clk), .Q(\mem[12][1] ) );
  DFQD1 \mem_reg[12][0]  ( .D(n4461), .CP(clk), .Q(\mem[12][0] ) );
  DFQD1 \mem_reg[13][15]  ( .D(n4460), .CP(clk), .Q(\mem[13][15] ) );
  DFQD1 \mem_reg[13][14]  ( .D(n4459), .CP(clk), .Q(\mem[13][14] ) );
  DFQD1 \mem_reg[13][13]  ( .D(n4458), .CP(clk), .Q(\mem[13][13] ) );
  DFQD1 \mem_reg[13][12]  ( .D(n4457), .CP(clk), .Q(\mem[13][12] ) );
  DFQD1 \mem_reg[13][11]  ( .D(n4456), .CP(clk), .Q(\mem[13][11] ) );
  DFQD1 \mem_reg[13][10]  ( .D(n4455), .CP(clk), .Q(\mem[13][10] ) );
  DFQD1 \mem_reg[13][9]  ( .D(n4454), .CP(clk), .Q(\mem[13][9] ) );
  DFQD1 \mem_reg[13][8]  ( .D(n4453), .CP(clk), .Q(\mem[13][8] ) );
  DFQD1 \mem_reg[13][7]  ( .D(n4452), .CP(clk), .Q(\mem[13][7] ) );
  DFQD1 \mem_reg[13][6]  ( .D(n4451), .CP(clk), .Q(\mem[13][6] ) );
  DFQD1 \mem_reg[13][5]  ( .D(n4450), .CP(clk), .Q(\mem[13][5] ) );
  DFQD1 \mem_reg[13][4]  ( .D(n4449), .CP(clk), .Q(\mem[13][4] ) );
  DFQD1 \mem_reg[13][3]  ( .D(n4448), .CP(clk), .Q(\mem[13][3] ) );
  DFQD1 \mem_reg[13][2]  ( .D(n4447), .CP(clk), .Q(\mem[13][2] ) );
  DFQD1 \mem_reg[13][1]  ( .D(n4446), .CP(clk), .Q(\mem[13][1] ) );
  DFQD1 \mem_reg[13][0]  ( .D(n4445), .CP(clk), .Q(\mem[13][0] ) );
  DFQD1 \mem_reg[14][15]  ( .D(n4444), .CP(clk), .Q(\mem[14][15] ) );
  DFQD1 \mem_reg[14][14]  ( .D(n4443), .CP(clk), .Q(\mem[14][14] ) );
  DFQD1 \mem_reg[14][13]  ( .D(n4442), .CP(clk), .Q(\mem[14][13] ) );
  DFQD1 \mem_reg[14][12]  ( .D(n4441), .CP(clk), .Q(\mem[14][12] ) );
  DFQD1 \mem_reg[14][11]  ( .D(n4440), .CP(clk), .Q(\mem[14][11] ) );
  DFQD1 \mem_reg[14][10]  ( .D(n4439), .CP(clk), .Q(\mem[14][10] ) );
  DFQD1 \mem_reg[14][9]  ( .D(n4438), .CP(clk), .Q(\mem[14][9] ) );
  DFQD1 \mem_reg[14][8]  ( .D(n4437), .CP(clk), .Q(\mem[14][8] ) );
  DFQD1 \mem_reg[14][7]  ( .D(n4436), .CP(clk), .Q(\mem[14][7] ) );
  DFQD1 \mem_reg[14][6]  ( .D(n4435), .CP(clk), .Q(\mem[14][6] ) );
  DFQD1 \mem_reg[14][5]  ( .D(n4434), .CP(clk), .Q(\mem[14][5] ) );
  DFQD1 \mem_reg[14][4]  ( .D(n4433), .CP(clk), .Q(\mem[14][4] ) );
  DFQD1 \mem_reg[14][3]  ( .D(n4432), .CP(clk), .Q(\mem[14][3] ) );
  DFQD1 \mem_reg[14][2]  ( .D(n4431), .CP(clk), .Q(\mem[14][2] ) );
  DFQD1 \mem_reg[14][1]  ( .D(n4430), .CP(clk), .Q(\mem[14][1] ) );
  DFQD1 \mem_reg[14][0]  ( .D(n4429), .CP(clk), .Q(\mem[14][0] ) );
  DFQD1 \mem_reg[15][15]  ( .D(n4428), .CP(clk), .Q(\mem[15][15] ) );
  DFQD1 \mem_reg[15][14]  ( .D(n4427), .CP(clk), .Q(\mem[15][14] ) );
  DFQD1 \mem_reg[15][13]  ( .D(n4426), .CP(clk), .Q(\mem[15][13] ) );
  DFQD1 \mem_reg[15][12]  ( .D(n4425), .CP(clk), .Q(\mem[15][12] ) );
  DFQD1 \mem_reg[15][11]  ( .D(n4424), .CP(clk), .Q(\mem[15][11] ) );
  DFQD1 \mem_reg[15][10]  ( .D(n4423), .CP(clk), .Q(\mem[15][10] ) );
  DFQD1 \mem_reg[15][9]  ( .D(n4422), .CP(clk), .Q(\mem[15][9] ) );
  DFQD1 \mem_reg[15][8]  ( .D(n4421), .CP(clk), .Q(\mem[15][8] ) );
  DFQD1 \mem_reg[15][7]  ( .D(n4420), .CP(clk), .Q(\mem[15][7] ) );
  DFQD1 \mem_reg[15][6]  ( .D(n4419), .CP(clk), .Q(\mem[15][6] ) );
  DFQD1 \mem_reg[15][5]  ( .D(n4418), .CP(clk), .Q(\mem[15][5] ) );
  DFQD1 \mem_reg[15][4]  ( .D(n4417), .CP(clk), .Q(\mem[15][4] ) );
  DFQD1 \mem_reg[15][3]  ( .D(n4416), .CP(clk), .Q(\mem[15][3] ) );
  DFQD1 \mem_reg[15][2]  ( .D(n4415), .CP(clk), .Q(\mem[15][2] ) );
  DFQD1 \mem_reg[15][1]  ( .D(n4414), .CP(clk), .Q(\mem[15][1] ) );
  DFQD1 \mem_reg[15][0]  ( .D(n4413), .CP(clk), .Q(\mem[15][0] ) );
  DFQD1 \mem_reg[16][15]  ( .D(n4412), .CP(clk), .Q(\mem[16][15] ) );
  DFQD1 \mem_reg[16][14]  ( .D(n4411), .CP(clk), .Q(\mem[16][14] ) );
  DFQD1 \mem_reg[16][13]  ( .D(n4410), .CP(clk), .Q(\mem[16][13] ) );
  DFQD1 \mem_reg[16][12]  ( .D(n4409), .CP(clk), .Q(\mem[16][12] ) );
  DFQD1 \mem_reg[16][11]  ( .D(n4408), .CP(clk), .Q(\mem[16][11] ) );
  DFQD1 \mem_reg[16][10]  ( .D(n4407), .CP(clk), .Q(\mem[16][10] ) );
  DFQD1 \mem_reg[16][9]  ( .D(n4406), .CP(clk), .Q(\mem[16][9] ) );
  DFQD1 \mem_reg[16][8]  ( .D(n4405), .CP(clk), .Q(\mem[16][8] ) );
  DFQD1 \mem_reg[16][7]  ( .D(n4404), .CP(clk), .Q(\mem[16][7] ) );
  DFQD1 \mem_reg[16][6]  ( .D(n4403), .CP(clk), .Q(\mem[16][6] ) );
  DFQD1 \mem_reg[16][5]  ( .D(n4402), .CP(clk), .Q(\mem[16][5] ) );
  DFQD1 \mem_reg[16][4]  ( .D(n4401), .CP(clk), .Q(\mem[16][4] ) );
  DFQD1 \mem_reg[16][3]  ( .D(n4400), .CP(clk), .Q(\mem[16][3] ) );
  DFQD1 \mem_reg[16][2]  ( .D(n4399), .CP(clk), .Q(\mem[16][2] ) );
  DFQD1 \mem_reg[16][1]  ( .D(n4398), .CP(clk), .Q(\mem[16][1] ) );
  DFQD1 \mem_reg[16][0]  ( .D(n4397), .CP(clk), .Q(\mem[16][0] ) );
  DFQD1 \mem_reg[17][15]  ( .D(n4396), .CP(clk), .Q(\mem[17][15] ) );
  DFQD1 \mem_reg[17][14]  ( .D(n4395), .CP(clk), .Q(\mem[17][14] ) );
  DFQD1 \mem_reg[17][13]  ( .D(n4394), .CP(clk), .Q(\mem[17][13] ) );
  DFQD1 \mem_reg[17][12]  ( .D(n4393), .CP(clk), .Q(\mem[17][12] ) );
  DFQD1 \mem_reg[17][11]  ( .D(n4392), .CP(clk), .Q(\mem[17][11] ) );
  DFQD1 \mem_reg[17][10]  ( .D(n4391), .CP(clk), .Q(\mem[17][10] ) );
  DFQD1 \mem_reg[17][9]  ( .D(n4390), .CP(clk), .Q(\mem[17][9] ) );
  DFQD1 \mem_reg[17][8]  ( .D(n4389), .CP(clk), .Q(\mem[17][8] ) );
  DFQD1 \mem_reg[17][7]  ( .D(n4388), .CP(clk), .Q(\mem[17][7] ) );
  DFQD1 \mem_reg[17][6]  ( .D(n4387), .CP(clk), .Q(\mem[17][6] ) );
  DFQD1 \mem_reg[17][5]  ( .D(n4386), .CP(clk), .Q(\mem[17][5] ) );
  DFQD1 \mem_reg[17][4]  ( .D(n4385), .CP(clk), .Q(\mem[17][4] ) );
  DFQD1 \mem_reg[17][3]  ( .D(n4384), .CP(clk), .Q(\mem[17][3] ) );
  DFQD1 \mem_reg[17][2]  ( .D(n4383), .CP(clk), .Q(\mem[17][2] ) );
  DFQD1 \mem_reg[17][1]  ( .D(n4382), .CP(clk), .Q(\mem[17][1] ) );
  DFQD1 \mem_reg[17][0]  ( .D(n4381), .CP(clk), .Q(\mem[17][0] ) );
  DFQD1 \mem_reg[18][15]  ( .D(n4380), .CP(clk), .Q(\mem[18][15] ) );
  DFQD1 \mem_reg[18][14]  ( .D(n4379), .CP(clk), .Q(\mem[18][14] ) );
  DFQD1 \mem_reg[18][13]  ( .D(n4378), .CP(clk), .Q(\mem[18][13] ) );
  DFQD1 \mem_reg[18][12]  ( .D(n4377), .CP(clk), .Q(\mem[18][12] ) );
  DFQD1 \mem_reg[18][11]  ( .D(n4376), .CP(clk), .Q(\mem[18][11] ) );
  DFQD1 \mem_reg[18][10]  ( .D(n4375), .CP(clk), .Q(\mem[18][10] ) );
  DFQD1 \mem_reg[18][9]  ( .D(n4374), .CP(clk), .Q(\mem[18][9] ) );
  DFQD1 \mem_reg[18][8]  ( .D(n4373), .CP(clk), .Q(\mem[18][8] ) );
  DFQD1 \mem_reg[18][7]  ( .D(n4372), .CP(clk), .Q(\mem[18][7] ) );
  DFQD1 \mem_reg[18][6]  ( .D(n4371), .CP(clk), .Q(\mem[18][6] ) );
  DFQD1 \mem_reg[18][5]  ( .D(n4370), .CP(clk), .Q(\mem[18][5] ) );
  DFQD1 \mem_reg[18][4]  ( .D(n4369), .CP(clk), .Q(\mem[18][4] ) );
  DFQD1 \mem_reg[18][3]  ( .D(n4368), .CP(clk), .Q(\mem[18][3] ) );
  DFQD1 \mem_reg[18][2]  ( .D(n4367), .CP(clk), .Q(\mem[18][2] ) );
  DFQD1 \mem_reg[18][1]  ( .D(n4366), .CP(clk), .Q(\mem[18][1] ) );
  DFQD1 \mem_reg[18][0]  ( .D(n4365), .CP(clk), .Q(\mem[18][0] ) );
  DFQD1 \mem_reg[19][15]  ( .D(n4364), .CP(clk), .Q(\mem[19][15] ) );
  DFQD1 \mem_reg[19][14]  ( .D(n4363), .CP(clk), .Q(\mem[19][14] ) );
  DFQD1 \mem_reg[19][13]  ( .D(n4362), .CP(clk), .Q(\mem[19][13] ) );
  DFQD1 \mem_reg[19][12]  ( .D(n4361), .CP(clk), .Q(\mem[19][12] ) );
  DFQD1 \mem_reg[19][11]  ( .D(n4360), .CP(clk), .Q(\mem[19][11] ) );
  DFQD1 \mem_reg[19][10]  ( .D(n4359), .CP(clk), .Q(\mem[19][10] ) );
  DFQD1 \mem_reg[19][9]  ( .D(n4358), .CP(clk), .Q(\mem[19][9] ) );
  DFQD1 \mem_reg[19][8]  ( .D(n4357), .CP(clk), .Q(\mem[19][8] ) );
  DFQD1 \mem_reg[19][7]  ( .D(n4356), .CP(clk), .Q(\mem[19][7] ) );
  DFQD1 \mem_reg[19][6]  ( .D(n4355), .CP(clk), .Q(\mem[19][6] ) );
  DFQD1 \mem_reg[19][5]  ( .D(n4354), .CP(clk), .Q(\mem[19][5] ) );
  DFQD1 \mem_reg[19][4]  ( .D(n4353), .CP(clk), .Q(\mem[19][4] ) );
  DFQD1 \mem_reg[19][3]  ( .D(n4352), .CP(clk), .Q(\mem[19][3] ) );
  DFQD1 \mem_reg[19][2]  ( .D(n4351), .CP(clk), .Q(\mem[19][2] ) );
  DFQD1 \mem_reg[19][1]  ( .D(n4350), .CP(clk), .Q(\mem[19][1] ) );
  DFQD1 \mem_reg[19][0]  ( .D(n4349), .CP(clk), .Q(\mem[19][0] ) );
  DFQD1 \mem_reg[20][15]  ( .D(n4348), .CP(clk), .Q(\mem[20][15] ) );
  DFQD1 \mem_reg[20][14]  ( .D(n4347), .CP(clk), .Q(\mem[20][14] ) );
  DFQD1 \mem_reg[20][13]  ( .D(n4346), .CP(clk), .Q(\mem[20][13] ) );
  DFQD1 \mem_reg[20][12]  ( .D(n4345), .CP(clk), .Q(\mem[20][12] ) );
  DFQD1 \mem_reg[20][11]  ( .D(n4344), .CP(clk), .Q(\mem[20][11] ) );
  DFQD1 \mem_reg[20][10]  ( .D(n4343), .CP(clk), .Q(\mem[20][10] ) );
  DFQD1 \mem_reg[20][9]  ( .D(n4342), .CP(clk), .Q(\mem[20][9] ) );
  DFQD1 \mem_reg[20][8]  ( .D(n4341), .CP(clk), .Q(\mem[20][8] ) );
  DFQD1 \mem_reg[20][7]  ( .D(n4340), .CP(clk), .Q(\mem[20][7] ) );
  DFQD1 \mem_reg[20][6]  ( .D(n4339), .CP(clk), .Q(\mem[20][6] ) );
  DFQD1 \mem_reg[20][5]  ( .D(n4338), .CP(clk), .Q(\mem[20][5] ) );
  DFQD1 \mem_reg[20][4]  ( .D(n4337), .CP(clk), .Q(\mem[20][4] ) );
  DFQD1 \mem_reg[20][3]  ( .D(n4336), .CP(clk), .Q(\mem[20][3] ) );
  DFQD1 \mem_reg[20][2]  ( .D(n4335), .CP(clk), .Q(\mem[20][2] ) );
  DFQD1 \mem_reg[20][1]  ( .D(n4334), .CP(clk), .Q(\mem[20][1] ) );
  DFQD1 \mem_reg[20][0]  ( .D(n4333), .CP(clk), .Q(\mem[20][0] ) );
  DFQD1 \mem_reg[21][15]  ( .D(n4332), .CP(clk), .Q(\mem[21][15] ) );
  DFQD1 \mem_reg[21][14]  ( .D(n4331), .CP(clk), .Q(\mem[21][14] ) );
  DFQD1 \mem_reg[21][13]  ( .D(n4330), .CP(clk), .Q(\mem[21][13] ) );
  DFQD1 \mem_reg[21][12]  ( .D(n4329), .CP(clk), .Q(\mem[21][12] ) );
  DFQD1 \mem_reg[21][11]  ( .D(n4328), .CP(clk), .Q(\mem[21][11] ) );
  DFQD1 \mem_reg[21][10]  ( .D(n4327), .CP(clk), .Q(\mem[21][10] ) );
  DFQD1 \mem_reg[21][9]  ( .D(n4326), .CP(clk), .Q(\mem[21][9] ) );
  DFQD1 \mem_reg[21][8]  ( .D(n4325), .CP(clk), .Q(\mem[21][8] ) );
  DFQD1 \mem_reg[21][7]  ( .D(n4324), .CP(clk), .Q(\mem[21][7] ) );
  DFQD1 \mem_reg[21][6]  ( .D(n4323), .CP(clk), .Q(\mem[21][6] ) );
  DFQD1 \mem_reg[21][5]  ( .D(n4322), .CP(clk), .Q(\mem[21][5] ) );
  DFQD1 \mem_reg[21][4]  ( .D(n4321), .CP(clk), .Q(\mem[21][4] ) );
  DFQD1 \mem_reg[21][3]  ( .D(n4320), .CP(clk), .Q(\mem[21][3] ) );
  DFQD1 \mem_reg[21][2]  ( .D(n4319), .CP(clk), .Q(\mem[21][2] ) );
  DFQD1 \mem_reg[21][1]  ( .D(n4318), .CP(clk), .Q(\mem[21][1] ) );
  DFQD1 \mem_reg[21][0]  ( .D(n4317), .CP(clk), .Q(\mem[21][0] ) );
  DFQD1 \mem_reg[22][15]  ( .D(n4316), .CP(clk), .Q(\mem[22][15] ) );
  DFQD1 \mem_reg[22][14]  ( .D(n4315), .CP(clk), .Q(\mem[22][14] ) );
  DFQD1 \mem_reg[22][13]  ( .D(n4314), .CP(clk), .Q(\mem[22][13] ) );
  DFQD1 \mem_reg[22][12]  ( .D(n4313), .CP(clk), .Q(\mem[22][12] ) );
  DFQD1 \mem_reg[22][11]  ( .D(n4312), .CP(clk), .Q(\mem[22][11] ) );
  DFQD1 \mem_reg[22][10]  ( .D(n4311), .CP(clk), .Q(\mem[22][10] ) );
  DFQD1 \mem_reg[22][9]  ( .D(n4310), .CP(clk), .Q(\mem[22][9] ) );
  DFQD1 \mem_reg[22][8]  ( .D(n4309), .CP(clk), .Q(\mem[22][8] ) );
  DFQD1 \mem_reg[22][7]  ( .D(n4308), .CP(clk), .Q(\mem[22][7] ) );
  DFQD1 \mem_reg[22][6]  ( .D(n4307), .CP(clk), .Q(\mem[22][6] ) );
  DFQD1 \mem_reg[22][5]  ( .D(n4306), .CP(clk), .Q(\mem[22][5] ) );
  DFQD1 \mem_reg[22][4]  ( .D(n4305), .CP(clk), .Q(\mem[22][4] ) );
  DFQD1 \mem_reg[22][3]  ( .D(n4304), .CP(clk), .Q(\mem[22][3] ) );
  DFQD1 \mem_reg[22][2]  ( .D(n4303), .CP(clk), .Q(\mem[22][2] ) );
  DFQD1 \mem_reg[22][1]  ( .D(n4302), .CP(clk), .Q(\mem[22][1] ) );
  DFQD1 \mem_reg[22][0]  ( .D(n4301), .CP(clk), .Q(\mem[22][0] ) );
  DFQD1 \mem_reg[23][15]  ( .D(n4300), .CP(clk), .Q(\mem[23][15] ) );
  DFQD1 \mem_reg[23][14]  ( .D(n4299), .CP(clk), .Q(\mem[23][14] ) );
  DFQD1 \mem_reg[23][13]  ( .D(n4298), .CP(clk), .Q(\mem[23][13] ) );
  DFQD1 \mem_reg[23][12]  ( .D(n4297), .CP(clk), .Q(\mem[23][12] ) );
  DFQD1 \mem_reg[23][11]  ( .D(n4296), .CP(clk), .Q(\mem[23][11] ) );
  DFQD1 \mem_reg[23][10]  ( .D(n4295), .CP(clk), .Q(\mem[23][10] ) );
  DFQD1 \mem_reg[23][9]  ( .D(n4294), .CP(clk), .Q(\mem[23][9] ) );
  DFQD1 \mem_reg[23][8]  ( .D(n4293), .CP(clk), .Q(\mem[23][8] ) );
  DFQD1 \mem_reg[23][7]  ( .D(n4292), .CP(clk), .Q(\mem[23][7] ) );
  DFQD1 \mem_reg[23][6]  ( .D(n4291), .CP(clk), .Q(\mem[23][6] ) );
  DFQD1 \mem_reg[23][5]  ( .D(n4290), .CP(clk), .Q(\mem[23][5] ) );
  DFQD1 \mem_reg[23][4]  ( .D(n4289), .CP(clk), .Q(\mem[23][4] ) );
  DFQD1 \mem_reg[23][3]  ( .D(n4288), .CP(clk), .Q(\mem[23][3] ) );
  DFQD1 \mem_reg[23][2]  ( .D(n4287), .CP(clk), .Q(\mem[23][2] ) );
  DFQD1 \mem_reg[23][1]  ( .D(n4286), .CP(clk), .Q(\mem[23][1] ) );
  DFQD1 \mem_reg[23][0]  ( .D(n4285), .CP(clk), .Q(\mem[23][0] ) );
  DFQD1 \mem_reg[24][15]  ( .D(n4284), .CP(clk), .Q(\mem[24][15] ) );
  DFQD1 \mem_reg[24][14]  ( .D(n4283), .CP(clk), .Q(\mem[24][14] ) );
  DFQD1 \mem_reg[24][13]  ( .D(n4282), .CP(clk), .Q(\mem[24][13] ) );
  DFQD1 \mem_reg[24][12]  ( .D(n4281), .CP(clk), .Q(\mem[24][12] ) );
  DFQD1 \mem_reg[24][11]  ( .D(n4280), .CP(clk), .Q(\mem[24][11] ) );
  DFQD1 \mem_reg[24][10]  ( .D(n4279), .CP(clk), .Q(\mem[24][10] ) );
  DFQD1 \mem_reg[24][9]  ( .D(n4278), .CP(clk), .Q(\mem[24][9] ) );
  DFQD1 \mem_reg[24][8]  ( .D(n4277), .CP(clk), .Q(\mem[24][8] ) );
  DFQD1 \mem_reg[24][7]  ( .D(n4276), .CP(clk), .Q(\mem[24][7] ) );
  DFQD1 \mem_reg[24][6]  ( .D(n4275), .CP(clk), .Q(\mem[24][6] ) );
  DFQD1 \mem_reg[24][5]  ( .D(n4274), .CP(clk), .Q(\mem[24][5] ) );
  DFQD1 \mem_reg[24][4]  ( .D(n4273), .CP(clk), .Q(\mem[24][4] ) );
  DFQD1 \mem_reg[24][3]  ( .D(n4272), .CP(clk), .Q(\mem[24][3] ) );
  DFQD1 \mem_reg[24][2]  ( .D(n4271), .CP(clk), .Q(\mem[24][2] ) );
  DFQD1 \mem_reg[24][1]  ( .D(n4270), .CP(clk), .Q(\mem[24][1] ) );
  DFQD1 \mem_reg[24][0]  ( .D(n4269), .CP(clk), .Q(\mem[24][0] ) );
  DFQD1 \mem_reg[25][15]  ( .D(n4268), .CP(clk), .Q(\mem[25][15] ) );
  DFQD1 \mem_reg[25][14]  ( .D(n4267), .CP(clk), .Q(\mem[25][14] ) );
  DFQD1 \mem_reg[25][13]  ( .D(n4266), .CP(clk), .Q(\mem[25][13] ) );
  DFQD1 \mem_reg[25][12]  ( .D(n4265), .CP(clk), .Q(\mem[25][12] ) );
  DFQD1 \mem_reg[25][11]  ( .D(n4264), .CP(clk), .Q(\mem[25][11] ) );
  DFQD1 \mem_reg[25][10]  ( .D(n4263), .CP(clk), .Q(\mem[25][10] ) );
  DFQD1 \mem_reg[25][9]  ( .D(n4262), .CP(clk), .Q(\mem[25][9] ) );
  DFQD1 \mem_reg[25][8]  ( .D(n4261), .CP(clk), .Q(\mem[25][8] ) );
  DFQD1 \mem_reg[25][7]  ( .D(n4260), .CP(clk), .Q(\mem[25][7] ) );
  DFQD1 \mem_reg[25][6]  ( .D(n4259), .CP(clk), .Q(\mem[25][6] ) );
  DFQD1 \mem_reg[25][5]  ( .D(n4258), .CP(clk), .Q(\mem[25][5] ) );
  DFQD1 \mem_reg[25][4]  ( .D(n4257), .CP(clk), .Q(\mem[25][4] ) );
  DFQD1 \mem_reg[25][3]  ( .D(n4256), .CP(clk), .Q(\mem[25][3] ) );
  DFQD1 \mem_reg[25][2]  ( .D(n4255), .CP(clk), .Q(\mem[25][2] ) );
  DFQD1 \mem_reg[25][1]  ( .D(n4254), .CP(clk), .Q(\mem[25][1] ) );
  DFQD1 \mem_reg[25][0]  ( .D(n4253), .CP(clk), .Q(\mem[25][0] ) );
  DFQD1 \mem_reg[26][15]  ( .D(n4252), .CP(clk), .Q(\mem[26][15] ) );
  DFQD1 \mem_reg[26][14]  ( .D(n4251), .CP(clk), .Q(\mem[26][14] ) );
  DFQD1 \mem_reg[26][13]  ( .D(n4250), .CP(clk), .Q(\mem[26][13] ) );
  DFQD1 \mem_reg[26][12]  ( .D(n4249), .CP(clk), .Q(\mem[26][12] ) );
  DFQD1 \mem_reg[26][11]  ( .D(n4248), .CP(clk), .Q(\mem[26][11] ) );
  DFQD1 \mem_reg[26][10]  ( .D(n4247), .CP(clk), .Q(\mem[26][10] ) );
  DFQD1 \mem_reg[26][9]  ( .D(n4246), .CP(clk), .Q(\mem[26][9] ) );
  DFQD1 \mem_reg[26][8]  ( .D(n4245), .CP(clk), .Q(\mem[26][8] ) );
  DFQD1 \mem_reg[26][7]  ( .D(n4244), .CP(clk), .Q(\mem[26][7] ) );
  DFQD1 \mem_reg[26][6]  ( .D(n4243), .CP(clk), .Q(\mem[26][6] ) );
  DFQD1 \mem_reg[26][5]  ( .D(n4242), .CP(clk), .Q(\mem[26][5] ) );
  DFQD1 \mem_reg[26][4]  ( .D(n4241), .CP(clk), .Q(\mem[26][4] ) );
  DFQD1 \mem_reg[26][3]  ( .D(n4240), .CP(clk), .Q(\mem[26][3] ) );
  DFQD1 \mem_reg[26][2]  ( .D(n4239), .CP(clk), .Q(\mem[26][2] ) );
  DFQD1 \mem_reg[26][1]  ( .D(n4238), .CP(clk), .Q(\mem[26][1] ) );
  DFQD1 \mem_reg[26][0]  ( .D(n4237), .CP(clk), .Q(\mem[26][0] ) );
  DFQD1 \mem_reg[27][15]  ( .D(n4236), .CP(clk), .Q(\mem[27][15] ) );
  DFQD1 \mem_reg[27][14]  ( .D(n4235), .CP(clk), .Q(\mem[27][14] ) );
  DFQD1 \mem_reg[27][13]  ( .D(n4234), .CP(clk), .Q(\mem[27][13] ) );
  DFQD1 \mem_reg[27][12]  ( .D(n4233), .CP(clk), .Q(\mem[27][12] ) );
  DFQD1 \mem_reg[27][11]  ( .D(n4232), .CP(clk), .Q(\mem[27][11] ) );
  DFQD1 \mem_reg[27][10]  ( .D(n4231), .CP(clk), .Q(\mem[27][10] ) );
  DFQD1 \mem_reg[27][9]  ( .D(n4230), .CP(clk), .Q(\mem[27][9] ) );
  DFQD1 \mem_reg[27][8]  ( .D(n4229), .CP(clk), .Q(\mem[27][8] ) );
  DFQD1 \mem_reg[27][7]  ( .D(n4228), .CP(clk), .Q(\mem[27][7] ) );
  DFQD1 \mem_reg[27][6]  ( .D(n4227), .CP(clk), .Q(\mem[27][6] ) );
  DFQD1 \mem_reg[27][5]  ( .D(n4226), .CP(clk), .Q(\mem[27][5] ) );
  DFQD1 \mem_reg[27][4]  ( .D(n4225), .CP(clk), .Q(\mem[27][4] ) );
  DFQD1 \mem_reg[27][3]  ( .D(n4224), .CP(clk), .Q(\mem[27][3] ) );
  DFQD1 \mem_reg[27][2]  ( .D(n4223), .CP(clk), .Q(\mem[27][2] ) );
  DFQD1 \mem_reg[27][1]  ( .D(n4222), .CP(clk), .Q(\mem[27][1] ) );
  DFQD1 \mem_reg[27][0]  ( .D(n4221), .CP(clk), .Q(\mem[27][0] ) );
  DFQD1 \mem_reg[28][15]  ( .D(n4220), .CP(clk), .Q(\mem[28][15] ) );
  DFQD1 \mem_reg[28][14]  ( .D(n4219), .CP(clk), .Q(\mem[28][14] ) );
  DFQD1 \mem_reg[28][13]  ( .D(n4218), .CP(clk), .Q(\mem[28][13] ) );
  DFQD1 \mem_reg[28][12]  ( .D(n4217), .CP(clk), .Q(\mem[28][12] ) );
  DFQD1 \mem_reg[28][11]  ( .D(n4216), .CP(clk), .Q(\mem[28][11] ) );
  DFQD1 \mem_reg[28][10]  ( .D(n4215), .CP(clk), .Q(\mem[28][10] ) );
  DFQD1 \mem_reg[28][9]  ( .D(n4214), .CP(clk), .Q(\mem[28][9] ) );
  DFQD1 \mem_reg[28][8]  ( .D(n4213), .CP(clk), .Q(\mem[28][8] ) );
  DFQD1 \mem_reg[28][7]  ( .D(n4212), .CP(clk), .Q(\mem[28][7] ) );
  DFQD1 \mem_reg[28][6]  ( .D(n4211), .CP(clk), .Q(\mem[28][6] ) );
  DFQD1 \mem_reg[28][5]  ( .D(n4210), .CP(clk), .Q(\mem[28][5] ) );
  DFQD1 \mem_reg[28][4]  ( .D(n4209), .CP(clk), .Q(\mem[28][4] ) );
  DFQD1 \mem_reg[28][3]  ( .D(n4208), .CP(clk), .Q(\mem[28][3] ) );
  DFQD1 \mem_reg[28][2]  ( .D(n4207), .CP(clk), .Q(\mem[28][2] ) );
  DFQD1 \mem_reg[28][1]  ( .D(n4206), .CP(clk), .Q(\mem[28][1] ) );
  DFQD1 \mem_reg[28][0]  ( .D(n4205), .CP(clk), .Q(\mem[28][0] ) );
  DFQD1 \mem_reg[29][15]  ( .D(n4204), .CP(clk), .Q(\mem[29][15] ) );
  DFQD1 \mem_reg[29][14]  ( .D(n4203), .CP(clk), .Q(\mem[29][14] ) );
  DFQD1 \mem_reg[29][13]  ( .D(n4202), .CP(clk), .Q(\mem[29][13] ) );
  DFQD1 \mem_reg[29][12]  ( .D(n4201), .CP(clk), .Q(\mem[29][12] ) );
  DFQD1 \mem_reg[29][11]  ( .D(n4200), .CP(clk), .Q(\mem[29][11] ) );
  DFQD1 \mem_reg[29][10]  ( .D(n4199), .CP(clk), .Q(\mem[29][10] ) );
  DFQD1 \mem_reg[29][9]  ( .D(n4198), .CP(clk), .Q(\mem[29][9] ) );
  DFQD1 \mem_reg[29][8]  ( .D(n4197), .CP(clk), .Q(\mem[29][8] ) );
  DFQD1 \mem_reg[29][7]  ( .D(n4196), .CP(clk), .Q(\mem[29][7] ) );
  DFQD1 \mem_reg[29][6]  ( .D(n4195), .CP(clk), .Q(\mem[29][6] ) );
  DFQD1 \mem_reg[29][5]  ( .D(n4194), .CP(clk), .Q(\mem[29][5] ) );
  DFQD1 \mem_reg[29][4]  ( .D(n4193), .CP(clk), .Q(\mem[29][4] ) );
  DFQD1 \mem_reg[29][3]  ( .D(n4192), .CP(clk), .Q(\mem[29][3] ) );
  DFQD1 \mem_reg[29][2]  ( .D(n4191), .CP(clk), .Q(\mem[29][2] ) );
  DFQD1 \mem_reg[29][1]  ( .D(n4190), .CP(clk), .Q(\mem[29][1] ) );
  DFQD1 \mem_reg[29][0]  ( .D(n4189), .CP(clk), .Q(\mem[29][0] ) );
  DFQD1 \mem_reg[30][15]  ( .D(n4188), .CP(clk), .Q(\mem[30][15] ) );
  DFQD1 \mem_reg[30][14]  ( .D(n4187), .CP(clk), .Q(\mem[30][14] ) );
  DFQD1 \mem_reg[30][13]  ( .D(n4186), .CP(clk), .Q(\mem[30][13] ) );
  DFQD1 \mem_reg[30][12]  ( .D(n4185), .CP(clk), .Q(\mem[30][12] ) );
  DFQD1 \mem_reg[30][11]  ( .D(n4184), .CP(clk), .Q(\mem[30][11] ) );
  DFQD1 \mem_reg[30][10]  ( .D(n4183), .CP(clk), .Q(\mem[30][10] ) );
  DFQD1 \mem_reg[30][9]  ( .D(n4182), .CP(clk), .Q(\mem[30][9] ) );
  DFQD1 \mem_reg[30][8]  ( .D(n4181), .CP(clk), .Q(\mem[30][8] ) );
  DFQD1 \mem_reg[30][7]  ( .D(n4180), .CP(clk), .Q(\mem[30][7] ) );
  DFQD1 \mem_reg[30][6]  ( .D(n4179), .CP(clk), .Q(\mem[30][6] ) );
  DFQD1 \mem_reg[30][5]  ( .D(n4178), .CP(clk), .Q(\mem[30][5] ) );
  DFQD1 \mem_reg[30][4]  ( .D(n4177), .CP(clk), .Q(\mem[30][4] ) );
  DFQD1 \mem_reg[30][3]  ( .D(n4176), .CP(clk), .Q(\mem[30][3] ) );
  DFQD1 \mem_reg[30][2]  ( .D(n4175), .CP(clk), .Q(\mem[30][2] ) );
  DFQD1 \mem_reg[30][1]  ( .D(n4174), .CP(clk), .Q(\mem[30][1] ) );
  DFQD1 \mem_reg[30][0]  ( .D(n4173), .CP(clk), .Q(\mem[30][0] ) );
  DFQD1 \mem_reg[31][15]  ( .D(n4172), .CP(clk), .Q(\mem[31][15] ) );
  DFQD1 \mem_reg[31][14]  ( .D(n4171), .CP(clk), .Q(\mem[31][14] ) );
  DFQD1 \mem_reg[31][13]  ( .D(n4170), .CP(clk), .Q(\mem[31][13] ) );
  DFQD1 \mem_reg[31][12]  ( .D(n4169), .CP(clk), .Q(\mem[31][12] ) );
  DFQD1 \mem_reg[31][11]  ( .D(n4168), .CP(clk), .Q(\mem[31][11] ) );
  DFQD1 \mem_reg[31][10]  ( .D(n4167), .CP(clk), .Q(\mem[31][10] ) );
  DFQD1 \mem_reg[31][9]  ( .D(n4166), .CP(clk), .Q(\mem[31][9] ) );
  DFQD1 \mem_reg[31][8]  ( .D(n4165), .CP(clk), .Q(\mem[31][8] ) );
  DFQD1 \mem_reg[31][7]  ( .D(n4164), .CP(clk), .Q(\mem[31][7] ) );
  DFQD1 \mem_reg[31][6]  ( .D(n4163), .CP(clk), .Q(\mem[31][6] ) );
  DFQD1 \mem_reg[31][5]  ( .D(n4162), .CP(clk), .Q(\mem[31][5] ) );
  DFQD1 \mem_reg[31][4]  ( .D(n4161), .CP(clk), .Q(\mem[31][4] ) );
  DFQD1 \mem_reg[31][3]  ( .D(n4160), .CP(clk), .Q(\mem[31][3] ) );
  DFQD1 \mem_reg[31][2]  ( .D(n4159), .CP(clk), .Q(\mem[31][2] ) );
  DFQD1 \mem_reg[31][1]  ( .D(n4158), .CP(clk), .Q(\mem[31][1] ) );
  DFQD1 \mem_reg[31][0]  ( .D(n4157), .CP(clk), .Q(\mem[31][0] ) );
  DFQD1 \mem_reg[32][15]  ( .D(n4156), .CP(clk), .Q(\mem[32][15] ) );
  DFQD1 \mem_reg[32][14]  ( .D(n4155), .CP(clk), .Q(\mem[32][14] ) );
  DFQD1 \mem_reg[32][13]  ( .D(n4154), .CP(clk), .Q(\mem[32][13] ) );
  DFQD1 \mem_reg[32][12]  ( .D(n4153), .CP(clk), .Q(\mem[32][12] ) );
  DFQD1 \mem_reg[32][11]  ( .D(n4152), .CP(clk), .Q(\mem[32][11] ) );
  DFQD1 \mem_reg[32][10]  ( .D(n4151), .CP(clk), .Q(\mem[32][10] ) );
  DFQD1 \mem_reg[32][9]  ( .D(n4150), .CP(clk), .Q(\mem[32][9] ) );
  DFQD1 \mem_reg[32][8]  ( .D(n4149), .CP(clk), .Q(\mem[32][8] ) );
  DFQD1 \mem_reg[32][7]  ( .D(n4148), .CP(clk), .Q(\mem[32][7] ) );
  DFQD1 \mem_reg[32][6]  ( .D(n4147), .CP(clk), .Q(\mem[32][6] ) );
  DFQD1 \mem_reg[32][5]  ( .D(n4146), .CP(clk), .Q(\mem[32][5] ) );
  DFQD1 \mem_reg[32][4]  ( .D(n4145), .CP(clk), .Q(\mem[32][4] ) );
  DFQD1 \mem_reg[32][3]  ( .D(n4144), .CP(clk), .Q(\mem[32][3] ) );
  DFQD1 \mem_reg[32][2]  ( .D(n4143), .CP(clk), .Q(\mem[32][2] ) );
  DFQD1 \mem_reg[32][1]  ( .D(n4142), .CP(clk), .Q(\mem[32][1] ) );
  DFQD1 \mem_reg[32][0]  ( .D(n4141), .CP(clk), .Q(\mem[32][0] ) );
  DFQD1 \mem_reg[33][15]  ( .D(n4140), .CP(clk), .Q(\mem[33][15] ) );
  DFQD1 \mem_reg[33][14]  ( .D(n4139), .CP(clk), .Q(\mem[33][14] ) );
  DFQD1 \mem_reg[33][13]  ( .D(n4138), .CP(clk), .Q(\mem[33][13] ) );
  DFQD1 \mem_reg[33][12]  ( .D(n4137), .CP(clk), .Q(\mem[33][12] ) );
  DFQD1 \mem_reg[33][11]  ( .D(n4136), .CP(clk), .Q(\mem[33][11] ) );
  DFQD1 \mem_reg[33][10]  ( .D(n4135), .CP(clk), .Q(\mem[33][10] ) );
  DFQD1 \mem_reg[33][9]  ( .D(n4134), .CP(clk), .Q(\mem[33][9] ) );
  DFQD1 \mem_reg[33][8]  ( .D(n4133), .CP(clk), .Q(\mem[33][8] ) );
  DFQD1 \mem_reg[33][7]  ( .D(n4132), .CP(clk), .Q(\mem[33][7] ) );
  DFQD1 \mem_reg[33][6]  ( .D(n4131), .CP(clk), .Q(\mem[33][6] ) );
  DFQD1 \mem_reg[33][5]  ( .D(n4130), .CP(clk), .Q(\mem[33][5] ) );
  DFQD1 \mem_reg[33][4]  ( .D(n4129), .CP(clk), .Q(\mem[33][4] ) );
  DFQD1 \mem_reg[33][3]  ( .D(n4128), .CP(clk), .Q(\mem[33][3] ) );
  DFQD1 \mem_reg[33][2]  ( .D(n4127), .CP(clk), .Q(\mem[33][2] ) );
  DFQD1 \mem_reg[33][1]  ( .D(n4126), .CP(clk), .Q(\mem[33][1] ) );
  DFQD1 \mem_reg[33][0]  ( .D(n4125), .CP(clk), .Q(\mem[33][0] ) );
  DFQD1 \mem_reg[34][15]  ( .D(n4124), .CP(clk), .Q(\mem[34][15] ) );
  DFQD1 \mem_reg[34][14]  ( .D(n4123), .CP(clk), .Q(\mem[34][14] ) );
  DFQD1 \mem_reg[34][13]  ( .D(n4122), .CP(clk), .Q(\mem[34][13] ) );
  DFQD1 \mem_reg[34][12]  ( .D(n4121), .CP(clk), .Q(\mem[34][12] ) );
  DFQD1 \mem_reg[34][11]  ( .D(n4120), .CP(clk), .Q(\mem[34][11] ) );
  DFQD1 \mem_reg[34][10]  ( .D(n4119), .CP(clk), .Q(\mem[34][10] ) );
  DFQD1 \mem_reg[34][9]  ( .D(n4118), .CP(clk), .Q(\mem[34][9] ) );
  DFQD1 \mem_reg[34][8]  ( .D(n4117), .CP(clk), .Q(\mem[34][8] ) );
  DFQD1 \mem_reg[34][7]  ( .D(n4116), .CP(clk), .Q(\mem[34][7] ) );
  DFQD1 \mem_reg[34][6]  ( .D(n4115), .CP(clk), .Q(\mem[34][6] ) );
  DFQD1 \mem_reg[34][5]  ( .D(n4114), .CP(clk), .Q(\mem[34][5] ) );
  DFQD1 \mem_reg[34][4]  ( .D(n4113), .CP(clk), .Q(\mem[34][4] ) );
  DFQD1 \mem_reg[34][3]  ( .D(n4112), .CP(clk), .Q(\mem[34][3] ) );
  DFQD1 \mem_reg[34][2]  ( .D(n4111), .CP(clk), .Q(\mem[34][2] ) );
  DFQD1 \mem_reg[34][1]  ( .D(n4110), .CP(clk), .Q(\mem[34][1] ) );
  DFQD1 \mem_reg[34][0]  ( .D(n4109), .CP(clk), .Q(\mem[34][0] ) );
  DFQD1 \mem_reg[35][15]  ( .D(n4108), .CP(clk), .Q(\mem[35][15] ) );
  DFQD1 \mem_reg[35][14]  ( .D(n4107), .CP(clk), .Q(\mem[35][14] ) );
  DFQD1 \mem_reg[35][13]  ( .D(n4106), .CP(clk), .Q(\mem[35][13] ) );
  DFQD1 \mem_reg[35][12]  ( .D(n4105), .CP(clk), .Q(\mem[35][12] ) );
  DFQD1 \mem_reg[35][11]  ( .D(n4104), .CP(clk), .Q(\mem[35][11] ) );
  DFQD1 \mem_reg[35][10]  ( .D(n4103), .CP(clk), .Q(\mem[35][10] ) );
  DFQD1 \mem_reg[35][9]  ( .D(n4102), .CP(clk), .Q(\mem[35][9] ) );
  DFQD1 \mem_reg[35][8]  ( .D(n4101), .CP(clk), .Q(\mem[35][8] ) );
  DFQD1 \mem_reg[35][7]  ( .D(n4100), .CP(clk), .Q(\mem[35][7] ) );
  DFQD1 \mem_reg[35][6]  ( .D(n4099), .CP(clk), .Q(\mem[35][6] ) );
  DFQD1 \mem_reg[35][5]  ( .D(n4098), .CP(clk), .Q(\mem[35][5] ) );
  DFQD1 \mem_reg[35][4]  ( .D(n4097), .CP(clk), .Q(\mem[35][4] ) );
  DFQD1 \mem_reg[35][3]  ( .D(n4096), .CP(clk), .Q(\mem[35][3] ) );
  DFQD1 \mem_reg[35][2]  ( .D(n4095), .CP(clk), .Q(\mem[35][2] ) );
  DFQD1 \mem_reg[35][1]  ( .D(n4094), .CP(clk), .Q(\mem[35][1] ) );
  DFQD1 \mem_reg[35][0]  ( .D(n4093), .CP(clk), .Q(\mem[35][0] ) );
  DFQD1 \mem_reg[36][15]  ( .D(n4092), .CP(clk), .Q(\mem[36][15] ) );
  DFQD1 \mem_reg[36][14]  ( .D(n4091), .CP(clk), .Q(\mem[36][14] ) );
  DFQD1 \mem_reg[36][13]  ( .D(n4090), .CP(clk), .Q(\mem[36][13] ) );
  DFQD1 \mem_reg[36][12]  ( .D(n4089), .CP(clk), .Q(\mem[36][12] ) );
  DFQD1 \mem_reg[36][11]  ( .D(n4088), .CP(clk), .Q(\mem[36][11] ) );
  DFQD1 \mem_reg[36][10]  ( .D(n4087), .CP(clk), .Q(\mem[36][10] ) );
  DFQD1 \mem_reg[36][9]  ( .D(n4086), .CP(clk), .Q(\mem[36][9] ) );
  DFQD1 \mem_reg[36][8]  ( .D(n4085), .CP(clk), .Q(\mem[36][8] ) );
  DFQD1 \mem_reg[36][7]  ( .D(n4084), .CP(clk), .Q(\mem[36][7] ) );
  DFQD1 \mem_reg[36][6]  ( .D(n4083), .CP(clk), .Q(\mem[36][6] ) );
  DFQD1 \mem_reg[36][5]  ( .D(n4082), .CP(clk), .Q(\mem[36][5] ) );
  DFQD1 \mem_reg[36][4]  ( .D(n4081), .CP(clk), .Q(\mem[36][4] ) );
  DFQD1 \mem_reg[36][3]  ( .D(n4080), .CP(clk), .Q(\mem[36][3] ) );
  DFQD1 \mem_reg[36][2]  ( .D(n4079), .CP(clk), .Q(\mem[36][2] ) );
  DFQD1 \mem_reg[36][1]  ( .D(n4078), .CP(clk), .Q(\mem[36][1] ) );
  DFQD1 \mem_reg[36][0]  ( .D(n4077), .CP(clk), .Q(\mem[36][0] ) );
  DFQD1 \mem_reg[37][15]  ( .D(n4076), .CP(clk), .Q(\mem[37][15] ) );
  DFQD1 \mem_reg[37][14]  ( .D(n4075), .CP(clk), .Q(\mem[37][14] ) );
  DFQD1 \mem_reg[37][13]  ( .D(n4074), .CP(clk), .Q(\mem[37][13] ) );
  DFQD1 \mem_reg[37][12]  ( .D(n4073), .CP(clk), .Q(\mem[37][12] ) );
  DFQD1 \mem_reg[37][11]  ( .D(n4072), .CP(clk), .Q(\mem[37][11] ) );
  DFQD1 \mem_reg[37][10]  ( .D(n4071), .CP(clk), .Q(\mem[37][10] ) );
  DFQD1 \mem_reg[37][9]  ( .D(n4070), .CP(clk), .Q(\mem[37][9] ) );
  DFQD1 \mem_reg[37][8]  ( .D(n4069), .CP(clk), .Q(\mem[37][8] ) );
  DFQD1 \mem_reg[37][7]  ( .D(n4068), .CP(clk), .Q(\mem[37][7] ) );
  DFQD1 \mem_reg[37][6]  ( .D(n4067), .CP(clk), .Q(\mem[37][6] ) );
  DFQD1 \mem_reg[37][5]  ( .D(n4066), .CP(clk), .Q(\mem[37][5] ) );
  DFQD1 \mem_reg[37][4]  ( .D(n4065), .CP(clk), .Q(\mem[37][4] ) );
  DFQD1 \mem_reg[37][3]  ( .D(n4064), .CP(clk), .Q(\mem[37][3] ) );
  DFQD1 \mem_reg[37][2]  ( .D(n4063), .CP(clk), .Q(\mem[37][2] ) );
  DFQD1 \mem_reg[37][1]  ( .D(n4062), .CP(clk), .Q(\mem[37][1] ) );
  DFQD1 \mem_reg[37][0]  ( .D(n4061), .CP(clk), .Q(\mem[37][0] ) );
  DFQD1 \mem_reg[38][15]  ( .D(n4060), .CP(clk), .Q(\mem[38][15] ) );
  DFQD1 \mem_reg[38][14]  ( .D(n4059), .CP(clk), .Q(\mem[38][14] ) );
  DFQD1 \mem_reg[38][13]  ( .D(n4058), .CP(clk), .Q(\mem[38][13] ) );
  DFQD1 \mem_reg[38][12]  ( .D(n4057), .CP(clk), .Q(\mem[38][12] ) );
  DFQD1 \mem_reg[38][11]  ( .D(n4056), .CP(clk), .Q(\mem[38][11] ) );
  DFQD1 \mem_reg[38][10]  ( .D(n4055), .CP(clk), .Q(\mem[38][10] ) );
  DFQD1 \mem_reg[38][9]  ( .D(n4054), .CP(clk), .Q(\mem[38][9] ) );
  DFQD1 \mem_reg[38][8]  ( .D(n4053), .CP(clk), .Q(\mem[38][8] ) );
  DFQD1 \mem_reg[38][7]  ( .D(n4052), .CP(clk), .Q(\mem[38][7] ) );
  DFQD1 \mem_reg[38][6]  ( .D(n4051), .CP(clk), .Q(\mem[38][6] ) );
  DFQD1 \mem_reg[38][5]  ( .D(n4050), .CP(clk), .Q(\mem[38][5] ) );
  DFQD1 \mem_reg[38][4]  ( .D(n4049), .CP(clk), .Q(\mem[38][4] ) );
  DFQD1 \mem_reg[38][3]  ( .D(n4048), .CP(clk), .Q(\mem[38][3] ) );
  DFQD1 \mem_reg[38][2]  ( .D(n4047), .CP(clk), .Q(\mem[38][2] ) );
  DFQD1 \mem_reg[38][1]  ( .D(n4046), .CP(clk), .Q(\mem[38][1] ) );
  DFQD1 \mem_reg[38][0]  ( .D(n4045), .CP(clk), .Q(\mem[38][0] ) );
  DFQD1 \mem_reg[39][15]  ( .D(n4044), .CP(clk), .Q(\mem[39][15] ) );
  DFQD1 \mem_reg[39][14]  ( .D(n4043), .CP(clk), .Q(\mem[39][14] ) );
  DFQD1 \mem_reg[39][13]  ( .D(n4042), .CP(clk), .Q(\mem[39][13] ) );
  DFQD1 \mem_reg[39][12]  ( .D(n4041), .CP(clk), .Q(\mem[39][12] ) );
  DFQD1 \mem_reg[39][11]  ( .D(n4040), .CP(clk), .Q(\mem[39][11] ) );
  DFQD1 \mem_reg[39][10]  ( .D(n4039), .CP(clk), .Q(\mem[39][10] ) );
  DFQD1 \mem_reg[39][9]  ( .D(n4038), .CP(clk), .Q(\mem[39][9] ) );
  DFQD1 \mem_reg[39][8]  ( .D(n4037), .CP(clk), .Q(\mem[39][8] ) );
  DFQD1 \mem_reg[39][7]  ( .D(n4036), .CP(clk), .Q(\mem[39][7] ) );
  DFQD1 \mem_reg[39][6]  ( .D(n4035), .CP(clk), .Q(\mem[39][6] ) );
  DFQD1 \mem_reg[39][5]  ( .D(n4034), .CP(clk), .Q(\mem[39][5] ) );
  DFQD1 \mem_reg[39][4]  ( .D(n4033), .CP(clk), .Q(\mem[39][4] ) );
  DFQD1 \mem_reg[39][3]  ( .D(n4032), .CP(clk), .Q(\mem[39][3] ) );
  DFQD1 \mem_reg[39][2]  ( .D(n4031), .CP(clk), .Q(\mem[39][2] ) );
  DFQD1 \mem_reg[39][1]  ( .D(n4030), .CP(clk), .Q(\mem[39][1] ) );
  DFQD1 \mem_reg[39][0]  ( .D(n4029), .CP(clk), .Q(\mem[39][0] ) );
  DFQD1 \mem_reg[40][15]  ( .D(n4028), .CP(clk), .Q(\mem[40][15] ) );
  DFQD1 \mem_reg[40][14]  ( .D(n4027), .CP(clk), .Q(\mem[40][14] ) );
  DFQD1 \mem_reg[40][13]  ( .D(n4026), .CP(clk), .Q(\mem[40][13] ) );
  DFQD1 \mem_reg[40][12]  ( .D(n4025), .CP(clk), .Q(\mem[40][12] ) );
  DFQD1 \mem_reg[40][11]  ( .D(n4024), .CP(clk), .Q(\mem[40][11] ) );
  DFQD1 \mem_reg[40][10]  ( .D(n4023), .CP(clk), .Q(\mem[40][10] ) );
  DFQD1 \mem_reg[40][9]  ( .D(n4022), .CP(clk), .Q(\mem[40][9] ) );
  DFQD1 \mem_reg[40][8]  ( .D(n4021), .CP(clk), .Q(\mem[40][8] ) );
  DFQD1 \mem_reg[40][7]  ( .D(n4020), .CP(clk), .Q(\mem[40][7] ) );
  DFQD1 \mem_reg[40][6]  ( .D(n4019), .CP(clk), .Q(\mem[40][6] ) );
  DFQD1 \mem_reg[40][5]  ( .D(n4018), .CP(clk), .Q(\mem[40][5] ) );
  DFQD1 \mem_reg[40][4]  ( .D(n4017), .CP(clk), .Q(\mem[40][4] ) );
  DFQD1 \mem_reg[40][3]  ( .D(n4016), .CP(clk), .Q(\mem[40][3] ) );
  DFQD1 \mem_reg[40][2]  ( .D(n4015), .CP(clk), .Q(\mem[40][2] ) );
  DFQD1 \mem_reg[40][1]  ( .D(n4014), .CP(clk), .Q(\mem[40][1] ) );
  DFQD1 \mem_reg[40][0]  ( .D(n4013), .CP(clk), .Q(\mem[40][0] ) );
  DFQD1 \mem_reg[41][15]  ( .D(n4012), .CP(clk), .Q(\mem[41][15] ) );
  DFQD1 \mem_reg[41][14]  ( .D(n4011), .CP(clk), .Q(\mem[41][14] ) );
  DFQD1 \mem_reg[41][13]  ( .D(n4010), .CP(clk), .Q(\mem[41][13] ) );
  DFQD1 \mem_reg[41][12]  ( .D(n4009), .CP(clk), .Q(\mem[41][12] ) );
  DFQD1 \mem_reg[41][11]  ( .D(n4008), .CP(clk), .Q(\mem[41][11] ) );
  DFQD1 \mem_reg[41][10]  ( .D(n4007), .CP(clk), .Q(\mem[41][10] ) );
  DFQD1 \mem_reg[41][9]  ( .D(n4006), .CP(clk), .Q(\mem[41][9] ) );
  DFQD1 \mem_reg[41][8]  ( .D(n4005), .CP(clk), .Q(\mem[41][8] ) );
  DFQD1 \mem_reg[41][7]  ( .D(n4004), .CP(clk), .Q(\mem[41][7] ) );
  DFQD1 \mem_reg[41][6]  ( .D(n4003), .CP(clk), .Q(\mem[41][6] ) );
  DFQD1 \mem_reg[41][5]  ( .D(n4002), .CP(clk), .Q(\mem[41][5] ) );
  DFQD1 \mem_reg[41][4]  ( .D(n4001), .CP(clk), .Q(\mem[41][4] ) );
  DFQD1 \mem_reg[41][3]  ( .D(n4000), .CP(clk), .Q(\mem[41][3] ) );
  DFQD1 \mem_reg[41][2]  ( .D(n3999), .CP(clk), .Q(\mem[41][2] ) );
  DFQD1 \mem_reg[41][1]  ( .D(n3998), .CP(clk), .Q(\mem[41][1] ) );
  DFQD1 \mem_reg[41][0]  ( .D(n3997), .CP(clk), .Q(\mem[41][0] ) );
  DFQD1 \mem_reg[42][15]  ( .D(n3996), .CP(clk), .Q(\mem[42][15] ) );
  DFQD1 \mem_reg[42][14]  ( .D(n3995), .CP(clk), .Q(\mem[42][14] ) );
  DFQD1 \mem_reg[42][13]  ( .D(n3994), .CP(clk), .Q(\mem[42][13] ) );
  DFQD1 \mem_reg[42][12]  ( .D(n3993), .CP(clk), .Q(\mem[42][12] ) );
  DFQD1 \mem_reg[42][11]  ( .D(n3992), .CP(clk), .Q(\mem[42][11] ) );
  DFQD1 \mem_reg[42][10]  ( .D(n3991), .CP(clk), .Q(\mem[42][10] ) );
  DFQD1 \mem_reg[42][9]  ( .D(n3990), .CP(clk), .Q(\mem[42][9] ) );
  DFQD1 \mem_reg[42][8]  ( .D(n3989), .CP(clk), .Q(\mem[42][8] ) );
  DFQD1 \mem_reg[42][7]  ( .D(n3988), .CP(clk), .Q(\mem[42][7] ) );
  DFQD1 \mem_reg[42][6]  ( .D(n3987), .CP(clk), .Q(\mem[42][6] ) );
  DFQD1 \mem_reg[42][5]  ( .D(n3986), .CP(clk), .Q(\mem[42][5] ) );
  DFQD1 \mem_reg[42][4]  ( .D(n3985), .CP(clk), .Q(\mem[42][4] ) );
  DFQD1 \mem_reg[42][3]  ( .D(n3984), .CP(clk), .Q(\mem[42][3] ) );
  DFQD1 \mem_reg[42][2]  ( .D(n3983), .CP(clk), .Q(\mem[42][2] ) );
  DFQD1 \mem_reg[42][1]  ( .D(n3982), .CP(clk), .Q(\mem[42][1] ) );
  DFQD1 \mem_reg[42][0]  ( .D(n3981), .CP(clk), .Q(\mem[42][0] ) );
  DFQD1 \mem_reg[43][15]  ( .D(n3980), .CP(clk), .Q(\mem[43][15] ) );
  DFQD1 \mem_reg[43][14]  ( .D(n3979), .CP(clk), .Q(\mem[43][14] ) );
  DFQD1 \mem_reg[43][13]  ( .D(n3978), .CP(clk), .Q(\mem[43][13] ) );
  DFQD1 \mem_reg[43][12]  ( .D(n3977), .CP(clk), .Q(\mem[43][12] ) );
  DFQD1 \mem_reg[43][11]  ( .D(n3976), .CP(clk), .Q(\mem[43][11] ) );
  DFQD1 \mem_reg[43][10]  ( .D(n3975), .CP(clk), .Q(\mem[43][10] ) );
  DFQD1 \mem_reg[43][9]  ( .D(n3974), .CP(clk), .Q(\mem[43][9] ) );
  DFQD1 \mem_reg[43][8]  ( .D(n3973), .CP(clk), .Q(\mem[43][8] ) );
  DFQD1 \mem_reg[43][7]  ( .D(n3972), .CP(clk), .Q(\mem[43][7] ) );
  DFQD1 \mem_reg[43][6]  ( .D(n3971), .CP(clk), .Q(\mem[43][6] ) );
  DFQD1 \mem_reg[43][5]  ( .D(n3970), .CP(clk), .Q(\mem[43][5] ) );
  DFQD1 \mem_reg[43][4]  ( .D(n3969), .CP(clk), .Q(\mem[43][4] ) );
  DFQD1 \mem_reg[43][3]  ( .D(n3968), .CP(clk), .Q(\mem[43][3] ) );
  DFQD1 \mem_reg[43][2]  ( .D(n3967), .CP(clk), .Q(\mem[43][2] ) );
  DFQD1 \mem_reg[43][1]  ( .D(n3966), .CP(clk), .Q(\mem[43][1] ) );
  DFQD1 \mem_reg[43][0]  ( .D(n3965), .CP(clk), .Q(\mem[43][0] ) );
  DFQD1 \mem_reg[44][15]  ( .D(n3964), .CP(clk), .Q(\mem[44][15] ) );
  DFQD1 \mem_reg[44][14]  ( .D(n3963), .CP(clk), .Q(\mem[44][14] ) );
  DFQD1 \mem_reg[44][13]  ( .D(n3962), .CP(clk), .Q(\mem[44][13] ) );
  DFQD1 \mem_reg[44][12]  ( .D(n3961), .CP(clk), .Q(\mem[44][12] ) );
  DFQD1 \mem_reg[44][11]  ( .D(n3960), .CP(clk), .Q(\mem[44][11] ) );
  DFQD1 \mem_reg[44][10]  ( .D(n3959), .CP(clk), .Q(\mem[44][10] ) );
  DFQD1 \mem_reg[44][9]  ( .D(n3958), .CP(clk), .Q(\mem[44][9] ) );
  DFQD1 \mem_reg[44][8]  ( .D(n3957), .CP(clk), .Q(\mem[44][8] ) );
  DFQD1 \mem_reg[44][7]  ( .D(n3956), .CP(clk), .Q(\mem[44][7] ) );
  DFQD1 \mem_reg[44][6]  ( .D(n3955), .CP(clk), .Q(\mem[44][6] ) );
  DFQD1 \mem_reg[44][5]  ( .D(n3954), .CP(clk), .Q(\mem[44][5] ) );
  DFQD1 \mem_reg[44][4]  ( .D(n3953), .CP(clk), .Q(\mem[44][4] ) );
  DFQD1 \mem_reg[44][3]  ( .D(n3952), .CP(clk), .Q(\mem[44][3] ) );
  DFQD1 \mem_reg[44][2]  ( .D(n3951), .CP(clk), .Q(\mem[44][2] ) );
  DFQD1 \mem_reg[44][1]  ( .D(n3950), .CP(clk), .Q(\mem[44][1] ) );
  DFQD1 \mem_reg[44][0]  ( .D(n3949), .CP(clk), .Q(\mem[44][0] ) );
  DFQD1 \mem_reg[45][15]  ( .D(n3948), .CP(clk), .Q(\mem[45][15] ) );
  DFQD1 \mem_reg[45][14]  ( .D(n3947), .CP(clk), .Q(\mem[45][14] ) );
  DFQD1 \mem_reg[45][13]  ( .D(n3946), .CP(clk), .Q(\mem[45][13] ) );
  DFQD1 \mem_reg[45][12]  ( .D(n3945), .CP(clk), .Q(\mem[45][12] ) );
  DFQD1 \mem_reg[45][11]  ( .D(n3944), .CP(clk), .Q(\mem[45][11] ) );
  DFQD1 \mem_reg[45][10]  ( .D(n3943), .CP(clk), .Q(\mem[45][10] ) );
  DFQD1 \mem_reg[45][9]  ( .D(n3942), .CP(clk), .Q(\mem[45][9] ) );
  DFQD1 \mem_reg[45][8]  ( .D(n3941), .CP(clk), .Q(\mem[45][8] ) );
  DFQD1 \mem_reg[45][7]  ( .D(n3940), .CP(clk), .Q(\mem[45][7] ) );
  DFQD1 \mem_reg[45][6]  ( .D(n3939), .CP(clk), .Q(\mem[45][6] ) );
  DFQD1 \mem_reg[45][5]  ( .D(n3938), .CP(clk), .Q(\mem[45][5] ) );
  DFQD1 \mem_reg[45][4]  ( .D(n3937), .CP(clk), .Q(\mem[45][4] ) );
  DFQD1 \mem_reg[45][3]  ( .D(n3936), .CP(clk), .Q(\mem[45][3] ) );
  DFQD1 \mem_reg[45][2]  ( .D(n3935), .CP(clk), .Q(\mem[45][2] ) );
  DFQD1 \mem_reg[45][1]  ( .D(n3934), .CP(clk), .Q(\mem[45][1] ) );
  DFQD1 \mem_reg[45][0]  ( .D(n3933), .CP(clk), .Q(\mem[45][0] ) );
  DFQD1 \mem_reg[46][15]  ( .D(n3932), .CP(clk), .Q(\mem[46][15] ) );
  DFQD1 \mem_reg[46][14]  ( .D(n3931), .CP(clk), .Q(\mem[46][14] ) );
  DFQD1 \mem_reg[46][13]  ( .D(n3930), .CP(clk), .Q(\mem[46][13] ) );
  DFQD1 \mem_reg[46][12]  ( .D(n3929), .CP(clk), .Q(\mem[46][12] ) );
  DFQD1 \mem_reg[46][11]  ( .D(n3928), .CP(clk), .Q(\mem[46][11] ) );
  DFQD1 \mem_reg[46][10]  ( .D(n3927), .CP(clk), .Q(\mem[46][10] ) );
  DFQD1 \mem_reg[46][9]  ( .D(n3926), .CP(clk), .Q(\mem[46][9] ) );
  DFQD1 \mem_reg[46][8]  ( .D(n3925), .CP(clk), .Q(\mem[46][8] ) );
  DFQD1 \mem_reg[46][7]  ( .D(n3924), .CP(clk), .Q(\mem[46][7] ) );
  DFQD1 \mem_reg[46][6]  ( .D(n3923), .CP(clk), .Q(\mem[46][6] ) );
  DFQD1 \mem_reg[46][5]  ( .D(n3922), .CP(clk), .Q(\mem[46][5] ) );
  DFQD1 \mem_reg[46][4]  ( .D(n3921), .CP(clk), .Q(\mem[46][4] ) );
  DFQD1 \mem_reg[46][3]  ( .D(n3920), .CP(clk), .Q(\mem[46][3] ) );
  DFQD1 \mem_reg[46][2]  ( .D(n3919), .CP(clk), .Q(\mem[46][2] ) );
  DFQD1 \mem_reg[46][1]  ( .D(n3918), .CP(clk), .Q(\mem[46][1] ) );
  DFQD1 \mem_reg[46][0]  ( .D(n3917), .CP(clk), .Q(\mem[46][0] ) );
  DFQD1 \mem_reg[47][15]  ( .D(n3916), .CP(clk), .Q(\mem[47][15] ) );
  DFQD1 \mem_reg[47][14]  ( .D(n3915), .CP(clk), .Q(\mem[47][14] ) );
  DFQD1 \mem_reg[47][13]  ( .D(n3914), .CP(clk), .Q(\mem[47][13] ) );
  DFQD1 \mem_reg[47][12]  ( .D(n3913), .CP(clk), .Q(\mem[47][12] ) );
  DFQD1 \mem_reg[47][11]  ( .D(n3912), .CP(clk), .Q(\mem[47][11] ) );
  DFQD1 \mem_reg[47][10]  ( .D(n3911), .CP(clk), .Q(\mem[47][10] ) );
  DFQD1 \mem_reg[47][9]  ( .D(n3910), .CP(clk), .Q(\mem[47][9] ) );
  DFQD1 \mem_reg[47][8]  ( .D(n3909), .CP(clk), .Q(\mem[47][8] ) );
  DFQD1 \mem_reg[47][7]  ( .D(n3908), .CP(clk), .Q(\mem[47][7] ) );
  DFQD1 \mem_reg[47][6]  ( .D(n3907), .CP(clk), .Q(\mem[47][6] ) );
  DFQD1 \mem_reg[47][5]  ( .D(n3906), .CP(clk), .Q(\mem[47][5] ) );
  DFQD1 \mem_reg[47][4]  ( .D(n3905), .CP(clk), .Q(\mem[47][4] ) );
  DFQD1 \mem_reg[47][3]  ( .D(n3904), .CP(clk), .Q(\mem[47][3] ) );
  DFQD1 \mem_reg[47][2]  ( .D(n3903), .CP(clk), .Q(\mem[47][2] ) );
  DFQD1 \mem_reg[47][1]  ( .D(n3902), .CP(clk), .Q(\mem[47][1] ) );
  DFQD1 \mem_reg[47][0]  ( .D(n3901), .CP(clk), .Q(\mem[47][0] ) );
  DFQD1 \mem_reg[48][15]  ( .D(n3900), .CP(clk), .Q(\mem[48][15] ) );
  DFQD1 \mem_reg[48][14]  ( .D(n3899), .CP(clk), .Q(\mem[48][14] ) );
  DFQD1 \mem_reg[48][13]  ( .D(n3898), .CP(clk), .Q(\mem[48][13] ) );
  DFQD1 \mem_reg[48][12]  ( .D(n3897), .CP(clk), .Q(\mem[48][12] ) );
  DFQD1 \mem_reg[48][11]  ( .D(n3896), .CP(clk), .Q(\mem[48][11] ) );
  DFQD1 \mem_reg[48][10]  ( .D(n3895), .CP(clk), .Q(\mem[48][10] ) );
  DFQD1 \mem_reg[48][9]  ( .D(n3894), .CP(clk), .Q(\mem[48][9] ) );
  DFQD1 \mem_reg[48][8]  ( .D(n3893), .CP(clk), .Q(\mem[48][8] ) );
  DFQD1 \mem_reg[48][7]  ( .D(n3892), .CP(clk), .Q(\mem[48][7] ) );
  DFQD1 \mem_reg[48][6]  ( .D(n3891), .CP(clk), .Q(\mem[48][6] ) );
  DFQD1 \mem_reg[48][5]  ( .D(n3890), .CP(clk), .Q(\mem[48][5] ) );
  DFQD1 \mem_reg[48][4]  ( .D(n3889), .CP(clk), .Q(\mem[48][4] ) );
  DFQD1 \mem_reg[48][3]  ( .D(n3888), .CP(clk), .Q(\mem[48][3] ) );
  DFQD1 \mem_reg[48][2]  ( .D(n3887), .CP(clk), .Q(\mem[48][2] ) );
  DFQD1 \mem_reg[48][1]  ( .D(n3886), .CP(clk), .Q(\mem[48][1] ) );
  DFQD1 \mem_reg[48][0]  ( .D(n3885), .CP(clk), .Q(\mem[48][0] ) );
  DFQD1 \mem_reg[49][15]  ( .D(n3884), .CP(clk), .Q(\mem[49][15] ) );
  DFQD1 \mem_reg[49][14]  ( .D(n3883), .CP(clk), .Q(\mem[49][14] ) );
  DFQD1 \mem_reg[49][13]  ( .D(n3882), .CP(clk), .Q(\mem[49][13] ) );
  DFQD1 \mem_reg[49][12]  ( .D(n3881), .CP(clk), .Q(\mem[49][12] ) );
  DFQD1 \mem_reg[49][11]  ( .D(n3880), .CP(clk), .Q(\mem[49][11] ) );
  DFQD1 \mem_reg[49][10]  ( .D(n3879), .CP(clk), .Q(\mem[49][10] ) );
  DFQD1 \mem_reg[49][9]  ( .D(n3878), .CP(clk), .Q(\mem[49][9] ) );
  DFQD1 \mem_reg[49][8]  ( .D(n3877), .CP(clk), .Q(\mem[49][8] ) );
  DFQD1 \mem_reg[49][7]  ( .D(n3876), .CP(clk), .Q(\mem[49][7] ) );
  DFQD1 \mem_reg[49][6]  ( .D(n3875), .CP(clk), .Q(\mem[49][6] ) );
  DFQD1 \mem_reg[49][5]  ( .D(n3874), .CP(clk), .Q(\mem[49][5] ) );
  DFQD1 \mem_reg[49][4]  ( .D(n3873), .CP(clk), .Q(\mem[49][4] ) );
  DFQD1 \mem_reg[49][3]  ( .D(n3872), .CP(clk), .Q(\mem[49][3] ) );
  DFQD1 \mem_reg[49][2]  ( .D(n3871), .CP(clk), .Q(\mem[49][2] ) );
  DFQD1 \mem_reg[49][1]  ( .D(n3870), .CP(clk), .Q(\mem[49][1] ) );
  DFQD1 \mem_reg[49][0]  ( .D(n3869), .CP(clk), .Q(\mem[49][0] ) );
  DFQD1 \mem_reg[50][15]  ( .D(n3868), .CP(clk), .Q(\mem[50][15] ) );
  DFQD1 \mem_reg[50][14]  ( .D(n3867), .CP(clk), .Q(\mem[50][14] ) );
  DFQD1 \mem_reg[50][13]  ( .D(n3866), .CP(clk), .Q(\mem[50][13] ) );
  DFQD1 \mem_reg[50][12]  ( .D(n3865), .CP(clk), .Q(\mem[50][12] ) );
  DFQD1 \mem_reg[50][11]  ( .D(n3864), .CP(clk), .Q(\mem[50][11] ) );
  DFQD1 \mem_reg[50][10]  ( .D(n3863), .CP(clk), .Q(\mem[50][10] ) );
  DFQD1 \mem_reg[50][9]  ( .D(n3862), .CP(clk), .Q(\mem[50][9] ) );
  DFQD1 \mem_reg[50][8]  ( .D(n3861), .CP(clk), .Q(\mem[50][8] ) );
  DFQD1 \mem_reg[50][7]  ( .D(n3860), .CP(clk), .Q(\mem[50][7] ) );
  DFQD1 \mem_reg[50][6]  ( .D(n3859), .CP(clk), .Q(\mem[50][6] ) );
  DFQD1 \mem_reg[50][5]  ( .D(n3858), .CP(clk), .Q(\mem[50][5] ) );
  DFQD1 \mem_reg[50][4]  ( .D(n3857), .CP(clk), .Q(\mem[50][4] ) );
  DFQD1 \mem_reg[50][3]  ( .D(n3856), .CP(clk), .Q(\mem[50][3] ) );
  DFQD1 \mem_reg[50][2]  ( .D(n3855), .CP(clk), .Q(\mem[50][2] ) );
  DFQD1 \mem_reg[50][1]  ( .D(n3854), .CP(clk), .Q(\mem[50][1] ) );
  DFQD1 \mem_reg[50][0]  ( .D(n3853), .CP(clk), .Q(\mem[50][0] ) );
  DFQD1 \mem_reg[51][15]  ( .D(n3852), .CP(clk), .Q(\mem[51][15] ) );
  DFQD1 \mem_reg[51][14]  ( .D(n3851), .CP(clk), .Q(\mem[51][14] ) );
  DFQD1 \mem_reg[51][13]  ( .D(n3850), .CP(clk), .Q(\mem[51][13] ) );
  DFQD1 \mem_reg[51][12]  ( .D(n3849), .CP(clk), .Q(\mem[51][12] ) );
  DFQD1 \mem_reg[51][11]  ( .D(n3848), .CP(clk), .Q(\mem[51][11] ) );
  DFQD1 \mem_reg[51][10]  ( .D(n3847), .CP(clk), .Q(\mem[51][10] ) );
  DFQD1 \mem_reg[51][9]  ( .D(n3846), .CP(clk), .Q(\mem[51][9] ) );
  DFQD1 \mem_reg[51][8]  ( .D(n3845), .CP(clk), .Q(\mem[51][8] ) );
  DFQD1 \mem_reg[51][7]  ( .D(n3844), .CP(clk), .Q(\mem[51][7] ) );
  DFQD1 \mem_reg[51][6]  ( .D(n3843), .CP(clk), .Q(\mem[51][6] ) );
  DFQD1 \mem_reg[51][5]  ( .D(n3842), .CP(clk), .Q(\mem[51][5] ) );
  DFQD1 \mem_reg[51][4]  ( .D(n3841), .CP(clk), .Q(\mem[51][4] ) );
  DFQD1 \mem_reg[51][3]  ( .D(n3840), .CP(clk), .Q(\mem[51][3] ) );
  DFQD1 \mem_reg[51][2]  ( .D(n3839), .CP(clk), .Q(\mem[51][2] ) );
  DFQD1 \mem_reg[51][1]  ( .D(n3838), .CP(clk), .Q(\mem[51][1] ) );
  DFQD1 \mem_reg[51][0]  ( .D(n3837), .CP(clk), .Q(\mem[51][0] ) );
  DFQD1 \mem_reg[52][15]  ( .D(n3836), .CP(clk), .Q(\mem[52][15] ) );
  DFQD1 \mem_reg[52][14]  ( .D(n3835), .CP(clk), .Q(\mem[52][14] ) );
  DFQD1 \mem_reg[52][13]  ( .D(n3834), .CP(clk), .Q(\mem[52][13] ) );
  DFQD1 \mem_reg[52][12]  ( .D(n3833), .CP(clk), .Q(\mem[52][12] ) );
  DFQD1 \mem_reg[52][11]  ( .D(n3832), .CP(clk), .Q(\mem[52][11] ) );
  DFQD1 \mem_reg[52][10]  ( .D(n3831), .CP(clk), .Q(\mem[52][10] ) );
  DFQD1 \mem_reg[52][9]  ( .D(n3830), .CP(clk), .Q(\mem[52][9] ) );
  DFQD1 \mem_reg[52][8]  ( .D(n3829), .CP(clk), .Q(\mem[52][8] ) );
  DFQD1 \mem_reg[52][7]  ( .D(n3828), .CP(clk), .Q(\mem[52][7] ) );
  DFQD1 \mem_reg[52][6]  ( .D(n3827), .CP(clk), .Q(\mem[52][6] ) );
  DFQD1 \mem_reg[52][5]  ( .D(n3826), .CP(clk), .Q(\mem[52][5] ) );
  DFQD1 \mem_reg[52][4]  ( .D(n3825), .CP(clk), .Q(\mem[52][4] ) );
  DFQD1 \mem_reg[52][3]  ( .D(n3824), .CP(clk), .Q(\mem[52][3] ) );
  DFQD1 \mem_reg[52][2]  ( .D(n3823), .CP(clk), .Q(\mem[52][2] ) );
  DFQD1 \mem_reg[52][1]  ( .D(n3822), .CP(clk), .Q(\mem[52][1] ) );
  DFQD1 \mem_reg[52][0]  ( .D(n3821), .CP(clk), .Q(\mem[52][0] ) );
  DFQD1 \mem_reg[53][15]  ( .D(n3820), .CP(clk), .Q(\mem[53][15] ) );
  DFQD1 \mem_reg[53][14]  ( .D(n3819), .CP(clk), .Q(\mem[53][14] ) );
  DFQD1 \mem_reg[53][13]  ( .D(n3818), .CP(clk), .Q(\mem[53][13] ) );
  DFQD1 \mem_reg[53][12]  ( .D(n3817), .CP(clk), .Q(\mem[53][12] ) );
  DFQD1 \mem_reg[53][11]  ( .D(n3816), .CP(clk), .Q(\mem[53][11] ) );
  DFQD1 \mem_reg[53][10]  ( .D(n3815), .CP(clk), .Q(\mem[53][10] ) );
  DFQD1 \mem_reg[53][9]  ( .D(n3814), .CP(clk), .Q(\mem[53][9] ) );
  DFQD1 \mem_reg[53][8]  ( .D(n3813), .CP(clk), .Q(\mem[53][8] ) );
  DFQD1 \mem_reg[53][7]  ( .D(n3812), .CP(clk), .Q(\mem[53][7] ) );
  DFQD1 \mem_reg[53][6]  ( .D(n3811), .CP(clk), .Q(\mem[53][6] ) );
  DFQD1 \mem_reg[53][5]  ( .D(n3810), .CP(clk), .Q(\mem[53][5] ) );
  DFQD1 \mem_reg[53][4]  ( .D(n3809), .CP(clk), .Q(\mem[53][4] ) );
  DFQD1 \mem_reg[53][3]  ( .D(n3808), .CP(clk), .Q(\mem[53][3] ) );
  DFQD1 \mem_reg[53][2]  ( .D(n3807), .CP(clk), .Q(\mem[53][2] ) );
  DFQD1 \mem_reg[53][1]  ( .D(n3806), .CP(clk), .Q(\mem[53][1] ) );
  DFQD1 \mem_reg[53][0]  ( .D(n3805), .CP(clk), .Q(\mem[53][0] ) );
  DFQD1 \mem_reg[54][15]  ( .D(n3804), .CP(clk), .Q(\mem[54][15] ) );
  DFQD1 \mem_reg[54][14]  ( .D(n3803), .CP(clk), .Q(\mem[54][14] ) );
  DFQD1 \mem_reg[54][13]  ( .D(n3802), .CP(clk), .Q(\mem[54][13] ) );
  DFQD1 \mem_reg[54][12]  ( .D(n3801), .CP(clk), .Q(\mem[54][12] ) );
  DFQD1 \mem_reg[54][11]  ( .D(n3800), .CP(clk), .Q(\mem[54][11] ) );
  DFQD1 \mem_reg[54][10]  ( .D(n3799), .CP(clk), .Q(\mem[54][10] ) );
  DFQD1 \mem_reg[54][9]  ( .D(n3798), .CP(clk), .Q(\mem[54][9] ) );
  DFQD1 \mem_reg[54][8]  ( .D(n3797), .CP(clk), .Q(\mem[54][8] ) );
  DFQD1 \mem_reg[54][7]  ( .D(n3796), .CP(clk), .Q(\mem[54][7] ) );
  DFQD1 \mem_reg[54][6]  ( .D(n3795), .CP(clk), .Q(\mem[54][6] ) );
  DFQD1 \mem_reg[54][5]  ( .D(n3794), .CP(clk), .Q(\mem[54][5] ) );
  DFQD1 \mem_reg[54][4]  ( .D(n3793), .CP(clk), .Q(\mem[54][4] ) );
  DFQD1 \mem_reg[54][3]  ( .D(n3792), .CP(clk), .Q(\mem[54][3] ) );
  DFQD1 \mem_reg[54][2]  ( .D(n3791), .CP(clk), .Q(\mem[54][2] ) );
  DFQD1 \mem_reg[54][1]  ( .D(n3790), .CP(clk), .Q(\mem[54][1] ) );
  DFQD1 \mem_reg[54][0]  ( .D(n3789), .CP(clk), .Q(\mem[54][0] ) );
  DFQD1 \mem_reg[55][15]  ( .D(n3788), .CP(clk), .Q(\mem[55][15] ) );
  DFQD1 \mem_reg[55][14]  ( .D(n3787), .CP(clk), .Q(\mem[55][14] ) );
  DFQD1 \mem_reg[55][13]  ( .D(n3786), .CP(clk), .Q(\mem[55][13] ) );
  DFQD1 \mem_reg[55][12]  ( .D(n3785), .CP(clk), .Q(\mem[55][12] ) );
  DFQD1 \mem_reg[55][11]  ( .D(n3784), .CP(clk), .Q(\mem[55][11] ) );
  DFQD1 \mem_reg[55][10]  ( .D(n3783), .CP(clk), .Q(\mem[55][10] ) );
  DFQD1 \mem_reg[55][9]  ( .D(n3782), .CP(clk), .Q(\mem[55][9] ) );
  DFQD1 \mem_reg[55][8]  ( .D(n3781), .CP(clk), .Q(\mem[55][8] ) );
  DFQD1 \mem_reg[55][7]  ( .D(n3780), .CP(clk), .Q(\mem[55][7] ) );
  DFQD1 \mem_reg[55][6]  ( .D(n3779), .CP(clk), .Q(\mem[55][6] ) );
  DFQD1 \mem_reg[55][5]  ( .D(n3778), .CP(clk), .Q(\mem[55][5] ) );
  DFQD1 \mem_reg[55][4]  ( .D(n3777), .CP(clk), .Q(\mem[55][4] ) );
  DFQD1 \mem_reg[55][3]  ( .D(n3776), .CP(clk), .Q(\mem[55][3] ) );
  DFQD1 \mem_reg[55][2]  ( .D(n3775), .CP(clk), .Q(\mem[55][2] ) );
  DFQD1 \mem_reg[55][1]  ( .D(n3774), .CP(clk), .Q(\mem[55][1] ) );
  DFQD1 \mem_reg[55][0]  ( .D(n3773), .CP(clk), .Q(\mem[55][0] ) );
  DFQD1 \mem_reg[56][15]  ( .D(n3772), .CP(clk), .Q(\mem[56][15] ) );
  DFQD1 \mem_reg[56][14]  ( .D(n3771), .CP(clk), .Q(\mem[56][14] ) );
  DFQD1 \mem_reg[56][13]  ( .D(n3770), .CP(clk), .Q(\mem[56][13] ) );
  DFQD1 \mem_reg[56][12]  ( .D(n3769), .CP(clk), .Q(\mem[56][12] ) );
  DFQD1 \mem_reg[56][11]  ( .D(n3768), .CP(clk), .Q(\mem[56][11] ) );
  DFQD1 \mem_reg[56][10]  ( .D(n3767), .CP(clk), .Q(\mem[56][10] ) );
  DFQD1 \mem_reg[56][9]  ( .D(n3766), .CP(clk), .Q(\mem[56][9] ) );
  DFQD1 \mem_reg[56][8]  ( .D(n3765), .CP(clk), .Q(\mem[56][8] ) );
  DFQD1 \mem_reg[56][7]  ( .D(n3764), .CP(clk), .Q(\mem[56][7] ) );
  DFQD1 \mem_reg[56][6]  ( .D(n3763), .CP(clk), .Q(\mem[56][6] ) );
  DFQD1 \mem_reg[56][5]  ( .D(n3762), .CP(clk), .Q(\mem[56][5] ) );
  DFQD1 \mem_reg[56][4]  ( .D(n3761), .CP(clk), .Q(\mem[56][4] ) );
  DFQD1 \mem_reg[56][3]  ( .D(n3760), .CP(clk), .Q(\mem[56][3] ) );
  DFQD1 \mem_reg[56][2]  ( .D(n3759), .CP(clk), .Q(\mem[56][2] ) );
  DFQD1 \mem_reg[56][1]  ( .D(n3758), .CP(clk), .Q(\mem[56][1] ) );
  DFQD1 \mem_reg[56][0]  ( .D(n3757), .CP(clk), .Q(\mem[56][0] ) );
  DFQD1 \mem_reg[57][15]  ( .D(n3756), .CP(clk), .Q(\mem[57][15] ) );
  DFQD1 \mem_reg[57][14]  ( .D(n3755), .CP(clk), .Q(\mem[57][14] ) );
  DFQD1 \mem_reg[57][13]  ( .D(n3754), .CP(clk), .Q(\mem[57][13] ) );
  DFQD1 \mem_reg[57][12]  ( .D(n3753), .CP(clk), .Q(\mem[57][12] ) );
  DFQD1 \mem_reg[57][11]  ( .D(n3752), .CP(clk), .Q(\mem[57][11] ) );
  DFQD1 \mem_reg[57][10]  ( .D(n3751), .CP(clk), .Q(\mem[57][10] ) );
  DFQD1 \mem_reg[57][9]  ( .D(n3750), .CP(clk), .Q(\mem[57][9] ) );
  DFQD1 \mem_reg[57][8]  ( .D(n3749), .CP(clk), .Q(\mem[57][8] ) );
  DFQD1 \mem_reg[57][7]  ( .D(n3748), .CP(clk), .Q(\mem[57][7] ) );
  DFQD1 \mem_reg[57][6]  ( .D(n3747), .CP(clk), .Q(\mem[57][6] ) );
  DFQD1 \mem_reg[57][5]  ( .D(n3746), .CP(clk), .Q(\mem[57][5] ) );
  DFQD1 \mem_reg[57][4]  ( .D(n3745), .CP(clk), .Q(\mem[57][4] ) );
  DFQD1 \mem_reg[57][3]  ( .D(n3744), .CP(clk), .Q(\mem[57][3] ) );
  DFQD1 \mem_reg[57][2]  ( .D(n3743), .CP(clk), .Q(\mem[57][2] ) );
  DFQD1 \mem_reg[57][1]  ( .D(n3742), .CP(clk), .Q(\mem[57][1] ) );
  DFQD1 \mem_reg[57][0]  ( .D(n3741), .CP(clk), .Q(\mem[57][0] ) );
  DFQD1 \mem_reg[58][15]  ( .D(n3740), .CP(clk), .Q(\mem[58][15] ) );
  DFQD1 \mem_reg[58][14]  ( .D(n3739), .CP(clk), .Q(\mem[58][14] ) );
  DFQD1 \mem_reg[58][13]  ( .D(n3738), .CP(clk), .Q(\mem[58][13] ) );
  DFQD1 \mem_reg[58][12]  ( .D(n3737), .CP(clk), .Q(\mem[58][12] ) );
  DFQD1 \mem_reg[58][11]  ( .D(n3736), .CP(clk), .Q(\mem[58][11] ) );
  DFQD1 \mem_reg[58][10]  ( .D(n3735), .CP(clk), .Q(\mem[58][10] ) );
  DFQD1 \mem_reg[58][9]  ( .D(n3734), .CP(clk), .Q(\mem[58][9] ) );
  DFQD1 \mem_reg[58][8]  ( .D(n3733), .CP(clk), .Q(\mem[58][8] ) );
  DFQD1 \mem_reg[58][7]  ( .D(n3732), .CP(clk), .Q(\mem[58][7] ) );
  DFQD1 \mem_reg[58][6]  ( .D(n3731), .CP(clk), .Q(\mem[58][6] ) );
  DFQD1 \mem_reg[58][5]  ( .D(n3730), .CP(clk), .Q(\mem[58][5] ) );
  DFQD1 \mem_reg[58][4]  ( .D(n3729), .CP(clk), .Q(\mem[58][4] ) );
  DFQD1 \mem_reg[58][3]  ( .D(n3728), .CP(clk), .Q(\mem[58][3] ) );
  DFQD1 \mem_reg[58][2]  ( .D(n3727), .CP(clk), .Q(\mem[58][2] ) );
  DFQD1 \mem_reg[58][1]  ( .D(n3726), .CP(clk), .Q(\mem[58][1] ) );
  DFQD1 \mem_reg[58][0]  ( .D(n3725), .CP(clk), .Q(\mem[58][0] ) );
  DFQD1 \mem_reg[59][15]  ( .D(n3724), .CP(clk), .Q(\mem[59][15] ) );
  DFQD1 \mem_reg[59][14]  ( .D(n3723), .CP(clk), .Q(\mem[59][14] ) );
  DFQD1 \mem_reg[59][13]  ( .D(n3722), .CP(clk), .Q(\mem[59][13] ) );
  DFQD1 \mem_reg[59][12]  ( .D(n3721), .CP(clk), .Q(\mem[59][12] ) );
  DFQD1 \mem_reg[59][11]  ( .D(n3720), .CP(clk), .Q(\mem[59][11] ) );
  DFQD1 \mem_reg[59][10]  ( .D(n3719), .CP(clk), .Q(\mem[59][10] ) );
  DFQD1 \mem_reg[59][9]  ( .D(n3718), .CP(clk), .Q(\mem[59][9] ) );
  DFQD1 \mem_reg[59][8]  ( .D(n3717), .CP(clk), .Q(\mem[59][8] ) );
  DFQD1 \mem_reg[59][7]  ( .D(n3716), .CP(clk), .Q(\mem[59][7] ) );
  DFQD1 \mem_reg[59][6]  ( .D(n3715), .CP(clk), .Q(\mem[59][6] ) );
  DFQD1 \mem_reg[59][5]  ( .D(n3714), .CP(clk), .Q(\mem[59][5] ) );
  DFQD1 \mem_reg[59][4]  ( .D(n3713), .CP(clk), .Q(\mem[59][4] ) );
  DFQD1 \mem_reg[59][3]  ( .D(n3712), .CP(clk), .Q(\mem[59][3] ) );
  DFQD1 \mem_reg[59][2]  ( .D(n3711), .CP(clk), .Q(\mem[59][2] ) );
  DFQD1 \mem_reg[59][1]  ( .D(n3710), .CP(clk), .Q(\mem[59][1] ) );
  DFQD1 \mem_reg[59][0]  ( .D(n3709), .CP(clk), .Q(\mem[59][0] ) );
  DFQD1 \mem_reg[60][15]  ( .D(n3708), .CP(clk), .Q(\mem[60][15] ) );
  DFQD1 \mem_reg[60][14]  ( .D(n3707), .CP(clk), .Q(\mem[60][14] ) );
  DFQD1 \mem_reg[60][13]  ( .D(n3706), .CP(clk), .Q(\mem[60][13] ) );
  DFQD1 \mem_reg[60][12]  ( .D(n3705), .CP(clk), .Q(\mem[60][12] ) );
  DFQD1 \mem_reg[60][11]  ( .D(n3704), .CP(clk), .Q(\mem[60][11] ) );
  DFQD1 \mem_reg[60][10]  ( .D(n3703), .CP(clk), .Q(\mem[60][10] ) );
  DFQD1 \mem_reg[60][9]  ( .D(n3702), .CP(clk), .Q(\mem[60][9] ) );
  DFQD1 \mem_reg[60][8]  ( .D(n3701), .CP(clk), .Q(\mem[60][8] ) );
  DFQD1 \mem_reg[60][7]  ( .D(n3700), .CP(clk), .Q(\mem[60][7] ) );
  DFQD1 \mem_reg[60][6]  ( .D(n3699), .CP(clk), .Q(\mem[60][6] ) );
  DFQD1 \mem_reg[60][5]  ( .D(n3698), .CP(clk), .Q(\mem[60][5] ) );
  DFQD1 \mem_reg[60][4]  ( .D(n3697), .CP(clk), .Q(\mem[60][4] ) );
  DFQD1 \mem_reg[60][3]  ( .D(n3696), .CP(clk), .Q(\mem[60][3] ) );
  DFQD1 \mem_reg[60][2]  ( .D(n3695), .CP(clk), .Q(\mem[60][2] ) );
  DFQD1 \mem_reg[60][1]  ( .D(n3694), .CP(clk), .Q(\mem[60][1] ) );
  DFQD1 \mem_reg[60][0]  ( .D(n3693), .CP(clk), .Q(\mem[60][0] ) );
  DFQD1 \mem_reg[61][15]  ( .D(n3692), .CP(clk), .Q(\mem[61][15] ) );
  DFQD1 \mem_reg[61][14]  ( .D(n3691), .CP(clk), .Q(\mem[61][14] ) );
  DFQD1 \mem_reg[61][13]  ( .D(n3690), .CP(clk), .Q(\mem[61][13] ) );
  DFQD1 \mem_reg[61][12]  ( .D(n3689), .CP(clk), .Q(\mem[61][12] ) );
  DFQD1 \mem_reg[61][11]  ( .D(n3688), .CP(clk), .Q(\mem[61][11] ) );
  DFQD1 \mem_reg[61][10]  ( .D(n3687), .CP(clk), .Q(\mem[61][10] ) );
  DFQD1 \mem_reg[61][9]  ( .D(n3686), .CP(clk), .Q(\mem[61][9] ) );
  DFQD1 \mem_reg[61][8]  ( .D(n3685), .CP(clk), .Q(\mem[61][8] ) );
  DFQD1 \mem_reg[61][7]  ( .D(n3684), .CP(clk), .Q(\mem[61][7] ) );
  DFQD1 \mem_reg[61][6]  ( .D(n3683), .CP(clk), .Q(\mem[61][6] ) );
  DFQD1 \mem_reg[61][5]  ( .D(n3682), .CP(clk), .Q(\mem[61][5] ) );
  DFQD1 \mem_reg[61][4]  ( .D(n3681), .CP(clk), .Q(\mem[61][4] ) );
  DFQD1 \mem_reg[61][3]  ( .D(n3680), .CP(clk), .Q(\mem[61][3] ) );
  DFQD1 \mem_reg[61][2]  ( .D(n3679), .CP(clk), .Q(\mem[61][2] ) );
  DFQD1 \mem_reg[61][1]  ( .D(n3678), .CP(clk), .Q(\mem[61][1] ) );
  DFQD1 \mem_reg[61][0]  ( .D(n3677), .CP(clk), .Q(\mem[61][0] ) );
  DFQD1 \mem_reg[62][15]  ( .D(n3676), .CP(clk), .Q(\mem[62][15] ) );
  DFQD1 \mem_reg[62][14]  ( .D(n3675), .CP(clk), .Q(\mem[62][14] ) );
  DFQD1 \mem_reg[62][13]  ( .D(n3674), .CP(clk), .Q(\mem[62][13] ) );
  DFQD1 \mem_reg[62][12]  ( .D(n3673), .CP(clk), .Q(\mem[62][12] ) );
  DFQD1 \mem_reg[62][11]  ( .D(n3672), .CP(clk), .Q(\mem[62][11] ) );
  DFQD1 \mem_reg[62][10]  ( .D(n3671), .CP(clk), .Q(\mem[62][10] ) );
  DFQD1 \mem_reg[62][9]  ( .D(n3670), .CP(clk), .Q(\mem[62][9] ) );
  DFQD1 \mem_reg[62][8]  ( .D(n3669), .CP(clk), .Q(\mem[62][8] ) );
  DFQD1 \mem_reg[62][7]  ( .D(n3668), .CP(clk), .Q(\mem[62][7] ) );
  DFQD1 \mem_reg[62][6]  ( .D(n3667), .CP(clk), .Q(\mem[62][6] ) );
  DFQD1 \mem_reg[62][5]  ( .D(n3666), .CP(clk), .Q(\mem[62][5] ) );
  DFQD1 \mem_reg[62][4]  ( .D(n3665), .CP(clk), .Q(\mem[62][4] ) );
  DFQD1 \mem_reg[62][3]  ( .D(n3664), .CP(clk), .Q(\mem[62][3] ) );
  DFQD1 \mem_reg[62][2]  ( .D(n3663), .CP(clk), .Q(\mem[62][2] ) );
  DFQD1 \mem_reg[62][1]  ( .D(n3662), .CP(clk), .Q(\mem[62][1] ) );
  DFQD1 \mem_reg[62][0]  ( .D(n3661), .CP(clk), .Q(\mem[62][0] ) );
  DFQD1 \mem_reg[63][15]  ( .D(n3660), .CP(clk), .Q(\mem[63][15] ) );
  DFQD1 \mem_reg[63][14]  ( .D(n3659), .CP(clk), .Q(\mem[63][14] ) );
  DFQD1 \mem_reg[63][13]  ( .D(n3658), .CP(clk), .Q(\mem[63][13] ) );
  DFQD1 \mem_reg[63][12]  ( .D(n3657), .CP(clk), .Q(\mem[63][12] ) );
  DFQD1 \mem_reg[63][11]  ( .D(n3656), .CP(clk), .Q(\mem[63][11] ) );
  DFQD1 \mem_reg[63][10]  ( .D(n3655), .CP(clk), .Q(\mem[63][10] ) );
  DFQD1 \mem_reg[63][9]  ( .D(n3654), .CP(clk), .Q(\mem[63][9] ) );
  DFQD1 \mem_reg[63][8]  ( .D(n3653), .CP(clk), .Q(\mem[63][8] ) );
  DFQD1 \mem_reg[63][7]  ( .D(n3652), .CP(clk), .Q(\mem[63][7] ) );
  DFQD1 \mem_reg[63][6]  ( .D(n3651), .CP(clk), .Q(\mem[63][6] ) );
  DFQD1 \mem_reg[63][5]  ( .D(n3650), .CP(clk), .Q(\mem[63][5] ) );
  DFQD1 \mem_reg[63][4]  ( .D(n3649), .CP(clk), .Q(\mem[63][4] ) );
  DFQD1 \mem_reg[63][3]  ( .D(n3648), .CP(clk), .Q(\mem[63][3] ) );
  DFQD1 \mem_reg[63][2]  ( .D(n3647), .CP(clk), .Q(\mem[63][2] ) );
  DFQD1 \mem_reg[63][1]  ( .D(n3646), .CP(clk), .Q(\mem[63][1] ) );
  DFQD1 \mem_reg[63][0]  ( .D(n3645), .CP(clk), .Q(\mem[63][0] ) );
  DFQD1 \mem_reg[64][15]  ( .D(n3644), .CP(clk), .Q(\mem[64][15] ) );
  DFQD1 \mem_reg[64][14]  ( .D(n3643), .CP(clk), .Q(\mem[64][14] ) );
  DFQD1 \mem_reg[64][13]  ( .D(n3642), .CP(clk), .Q(\mem[64][13] ) );
  DFQD1 \mem_reg[64][12]  ( .D(n3641), .CP(clk), .Q(\mem[64][12] ) );
  DFQD1 \mem_reg[64][11]  ( .D(n3640), .CP(clk), .Q(\mem[64][11] ) );
  DFQD1 \mem_reg[64][10]  ( .D(n3639), .CP(clk), .Q(\mem[64][10] ) );
  DFQD1 \mem_reg[64][9]  ( .D(n3638), .CP(clk), .Q(\mem[64][9] ) );
  DFQD1 \mem_reg[64][8]  ( .D(n3637), .CP(clk), .Q(\mem[64][8] ) );
  DFQD1 \mem_reg[64][7]  ( .D(n3636), .CP(clk), .Q(\mem[64][7] ) );
  DFQD1 \mem_reg[64][6]  ( .D(n3635), .CP(clk), .Q(\mem[64][6] ) );
  DFQD1 \mem_reg[64][5]  ( .D(n3634), .CP(clk), .Q(\mem[64][5] ) );
  DFQD1 \mem_reg[64][4]  ( .D(n3633), .CP(clk), .Q(\mem[64][4] ) );
  DFQD1 \mem_reg[64][3]  ( .D(n3632), .CP(clk), .Q(\mem[64][3] ) );
  DFQD1 \mem_reg[64][2]  ( .D(n3631), .CP(clk), .Q(\mem[64][2] ) );
  DFQD1 \mem_reg[64][1]  ( .D(n3630), .CP(clk), .Q(\mem[64][1] ) );
  DFQD1 \mem_reg[64][0]  ( .D(n3629), .CP(clk), .Q(\mem[64][0] ) );
  DFQD1 \mem_reg[65][15]  ( .D(n3628), .CP(clk), .Q(\mem[65][15] ) );
  DFQD1 \mem_reg[65][14]  ( .D(n3627), .CP(clk), .Q(\mem[65][14] ) );
  DFQD1 \mem_reg[65][13]  ( .D(n3626), .CP(clk), .Q(\mem[65][13] ) );
  DFQD1 \mem_reg[65][12]  ( .D(n3625), .CP(clk), .Q(\mem[65][12] ) );
  DFQD1 \mem_reg[65][11]  ( .D(n3624), .CP(clk), .Q(\mem[65][11] ) );
  DFQD1 \mem_reg[65][10]  ( .D(n3623), .CP(clk), .Q(\mem[65][10] ) );
  DFQD1 \mem_reg[65][9]  ( .D(n3622), .CP(clk), .Q(\mem[65][9] ) );
  DFQD1 \mem_reg[65][8]  ( .D(n3621), .CP(clk), .Q(\mem[65][8] ) );
  DFQD1 \mem_reg[65][7]  ( .D(n3620), .CP(clk), .Q(\mem[65][7] ) );
  DFQD1 \mem_reg[65][6]  ( .D(n3619), .CP(clk), .Q(\mem[65][6] ) );
  DFQD1 \mem_reg[65][5]  ( .D(n3618), .CP(clk), .Q(\mem[65][5] ) );
  DFQD1 \mem_reg[65][4]  ( .D(n3617), .CP(clk), .Q(\mem[65][4] ) );
  DFQD1 \mem_reg[65][3]  ( .D(n3616), .CP(clk), .Q(\mem[65][3] ) );
  DFQD1 \mem_reg[65][2]  ( .D(n3615), .CP(clk), .Q(\mem[65][2] ) );
  DFQD1 \mem_reg[65][1]  ( .D(n3614), .CP(clk), .Q(\mem[65][1] ) );
  DFQD1 \mem_reg[65][0]  ( .D(n3613), .CP(clk), .Q(\mem[65][0] ) );
  DFQD1 \mem_reg[66][15]  ( .D(n3612), .CP(clk), .Q(\mem[66][15] ) );
  DFQD1 \mem_reg[66][14]  ( .D(n3611), .CP(clk), .Q(\mem[66][14] ) );
  DFQD1 \mem_reg[66][13]  ( .D(n3610), .CP(clk), .Q(\mem[66][13] ) );
  DFQD1 \mem_reg[66][12]  ( .D(n3609), .CP(clk), .Q(\mem[66][12] ) );
  DFQD1 \mem_reg[66][11]  ( .D(n3608), .CP(clk), .Q(\mem[66][11] ) );
  DFQD1 \mem_reg[66][10]  ( .D(n3607), .CP(clk), .Q(\mem[66][10] ) );
  DFQD1 \mem_reg[66][9]  ( .D(n3606), .CP(clk), .Q(\mem[66][9] ) );
  DFQD1 \mem_reg[66][8]  ( .D(n3605), .CP(clk), .Q(\mem[66][8] ) );
  DFQD1 \mem_reg[66][7]  ( .D(n3604), .CP(clk), .Q(\mem[66][7] ) );
  DFQD1 \mem_reg[66][6]  ( .D(n3603), .CP(clk), .Q(\mem[66][6] ) );
  DFQD1 \mem_reg[66][5]  ( .D(n3602), .CP(clk), .Q(\mem[66][5] ) );
  DFQD1 \mem_reg[66][4]  ( .D(n3601), .CP(clk), .Q(\mem[66][4] ) );
  DFQD1 \mem_reg[66][3]  ( .D(n3600), .CP(clk), .Q(\mem[66][3] ) );
  DFQD1 \mem_reg[66][2]  ( .D(n3599), .CP(clk), .Q(\mem[66][2] ) );
  DFQD1 \mem_reg[66][1]  ( .D(n3598), .CP(clk), .Q(\mem[66][1] ) );
  DFQD1 \mem_reg[66][0]  ( .D(n3597), .CP(clk), .Q(\mem[66][0] ) );
  DFQD1 \mem_reg[67][15]  ( .D(n3596), .CP(clk), .Q(\mem[67][15] ) );
  DFQD1 \mem_reg[67][14]  ( .D(n3595), .CP(clk), .Q(\mem[67][14] ) );
  DFQD1 \mem_reg[67][13]  ( .D(n3594), .CP(clk), .Q(\mem[67][13] ) );
  DFQD1 \mem_reg[67][12]  ( .D(n3593), .CP(clk), .Q(\mem[67][12] ) );
  DFQD1 \mem_reg[67][11]  ( .D(n3592), .CP(clk), .Q(\mem[67][11] ) );
  DFQD1 \mem_reg[67][10]  ( .D(n3591), .CP(clk), .Q(\mem[67][10] ) );
  DFQD1 \mem_reg[67][9]  ( .D(n3590), .CP(clk), .Q(\mem[67][9] ) );
  DFQD1 \mem_reg[67][8]  ( .D(n3589), .CP(clk), .Q(\mem[67][8] ) );
  DFQD1 \mem_reg[67][7]  ( .D(n3588), .CP(clk), .Q(\mem[67][7] ) );
  DFQD1 \mem_reg[67][6]  ( .D(n3587), .CP(clk), .Q(\mem[67][6] ) );
  DFQD1 \mem_reg[67][5]  ( .D(n3586), .CP(clk), .Q(\mem[67][5] ) );
  DFQD1 \mem_reg[67][4]  ( .D(n3585), .CP(clk), .Q(\mem[67][4] ) );
  DFQD1 \mem_reg[67][3]  ( .D(n3584), .CP(clk), .Q(\mem[67][3] ) );
  DFQD1 \mem_reg[67][2]  ( .D(n3583), .CP(clk), .Q(\mem[67][2] ) );
  DFQD1 \mem_reg[67][1]  ( .D(n3582), .CP(clk), .Q(\mem[67][1] ) );
  DFQD1 \mem_reg[67][0]  ( .D(n3581), .CP(clk), .Q(\mem[67][0] ) );
  DFQD1 \mem_reg[68][15]  ( .D(n3580), .CP(clk), .Q(\mem[68][15] ) );
  DFQD1 \mem_reg[68][14]  ( .D(n3579), .CP(clk), .Q(\mem[68][14] ) );
  DFQD1 \mem_reg[68][13]  ( .D(n3578), .CP(clk), .Q(\mem[68][13] ) );
  DFQD1 \mem_reg[68][12]  ( .D(n3577), .CP(clk), .Q(\mem[68][12] ) );
  DFQD1 \mem_reg[68][11]  ( .D(n3576), .CP(clk), .Q(\mem[68][11] ) );
  DFQD1 \mem_reg[68][10]  ( .D(n3575), .CP(clk), .Q(\mem[68][10] ) );
  DFQD1 \mem_reg[68][9]  ( .D(n3574), .CP(clk), .Q(\mem[68][9] ) );
  DFQD1 \mem_reg[68][8]  ( .D(n3573), .CP(clk), .Q(\mem[68][8] ) );
  DFQD1 \mem_reg[68][7]  ( .D(n3572), .CP(clk), .Q(\mem[68][7] ) );
  DFQD1 \mem_reg[68][6]  ( .D(n3571), .CP(clk), .Q(\mem[68][6] ) );
  DFQD1 \mem_reg[68][5]  ( .D(n3570), .CP(clk), .Q(\mem[68][5] ) );
  DFQD1 \mem_reg[68][4]  ( .D(n3569), .CP(clk), .Q(\mem[68][4] ) );
  DFQD1 \mem_reg[68][3]  ( .D(n3568), .CP(clk), .Q(\mem[68][3] ) );
  DFQD1 \mem_reg[68][2]  ( .D(n3567), .CP(clk), .Q(\mem[68][2] ) );
  DFQD1 \mem_reg[68][1]  ( .D(n3566), .CP(clk), .Q(\mem[68][1] ) );
  DFQD1 \mem_reg[68][0]  ( .D(n3565), .CP(clk), .Q(\mem[68][0] ) );
  DFQD1 \mem_reg[69][15]  ( .D(n3564), .CP(clk), .Q(\mem[69][15] ) );
  DFQD1 \mem_reg[69][14]  ( .D(n3563), .CP(clk), .Q(\mem[69][14] ) );
  DFQD1 \mem_reg[69][13]  ( .D(n3562), .CP(clk), .Q(\mem[69][13] ) );
  DFQD1 \mem_reg[69][12]  ( .D(n3561), .CP(clk), .Q(\mem[69][12] ) );
  DFQD1 \mem_reg[69][11]  ( .D(n3560), .CP(clk), .Q(\mem[69][11] ) );
  DFQD1 \mem_reg[69][10]  ( .D(n3559), .CP(clk), .Q(\mem[69][10] ) );
  DFQD1 \mem_reg[69][9]  ( .D(n3558), .CP(clk), .Q(\mem[69][9] ) );
  DFQD1 \mem_reg[69][8]  ( .D(n3557), .CP(clk), .Q(\mem[69][8] ) );
  DFQD1 \mem_reg[69][7]  ( .D(n3556), .CP(clk), .Q(\mem[69][7] ) );
  DFQD1 \mem_reg[69][6]  ( .D(n3555), .CP(clk), .Q(\mem[69][6] ) );
  DFQD1 \mem_reg[69][5]  ( .D(n3554), .CP(clk), .Q(\mem[69][5] ) );
  DFQD1 \mem_reg[69][4]  ( .D(n3553), .CP(clk), .Q(\mem[69][4] ) );
  DFQD1 \mem_reg[69][3]  ( .D(n3552), .CP(clk), .Q(\mem[69][3] ) );
  DFQD1 \mem_reg[69][2]  ( .D(n3551), .CP(clk), .Q(\mem[69][2] ) );
  DFQD1 \mem_reg[69][1]  ( .D(n3550), .CP(clk), .Q(\mem[69][1] ) );
  DFQD1 \mem_reg[69][0]  ( .D(n3549), .CP(clk), .Q(\mem[69][0] ) );
  DFQD1 \mem_reg[70][15]  ( .D(n3548), .CP(clk), .Q(\mem[70][15] ) );
  DFQD1 \mem_reg[70][14]  ( .D(n3547), .CP(clk), .Q(\mem[70][14] ) );
  DFQD1 \mem_reg[70][13]  ( .D(n3546), .CP(clk), .Q(\mem[70][13] ) );
  DFQD1 \mem_reg[70][12]  ( .D(n3545), .CP(clk), .Q(\mem[70][12] ) );
  DFQD1 \mem_reg[70][11]  ( .D(n3544), .CP(clk), .Q(\mem[70][11] ) );
  DFQD1 \mem_reg[70][10]  ( .D(n3543), .CP(clk), .Q(\mem[70][10] ) );
  DFQD1 \mem_reg[70][9]  ( .D(n3542), .CP(clk), .Q(\mem[70][9] ) );
  DFQD1 \mem_reg[70][8]  ( .D(n3541), .CP(clk), .Q(\mem[70][8] ) );
  DFQD1 \mem_reg[70][7]  ( .D(n3540), .CP(clk), .Q(\mem[70][7] ) );
  DFQD1 \mem_reg[70][6]  ( .D(n3539), .CP(clk), .Q(\mem[70][6] ) );
  DFQD1 \mem_reg[70][5]  ( .D(n3538), .CP(clk), .Q(\mem[70][5] ) );
  DFQD1 \mem_reg[70][4]  ( .D(n3537), .CP(clk), .Q(\mem[70][4] ) );
  DFQD1 \mem_reg[70][3]  ( .D(n3536), .CP(clk), .Q(\mem[70][3] ) );
  DFQD1 \mem_reg[70][2]  ( .D(n3535), .CP(clk), .Q(\mem[70][2] ) );
  DFQD1 \mem_reg[70][1]  ( .D(n3534), .CP(clk), .Q(\mem[70][1] ) );
  DFQD1 \mem_reg[70][0]  ( .D(n3533), .CP(clk), .Q(\mem[70][0] ) );
  DFQD1 \mem_reg[71][15]  ( .D(n3532), .CP(clk), .Q(\mem[71][15] ) );
  DFQD1 \mem_reg[71][14]  ( .D(n3531), .CP(clk), .Q(\mem[71][14] ) );
  DFQD1 \mem_reg[71][13]  ( .D(n3530), .CP(clk), .Q(\mem[71][13] ) );
  DFQD1 \mem_reg[71][12]  ( .D(n3529), .CP(clk), .Q(\mem[71][12] ) );
  DFQD1 \mem_reg[71][11]  ( .D(n3528), .CP(clk), .Q(\mem[71][11] ) );
  DFQD1 \mem_reg[71][10]  ( .D(n3527), .CP(clk), .Q(\mem[71][10] ) );
  DFQD1 \mem_reg[71][9]  ( .D(n3526), .CP(clk), .Q(\mem[71][9] ) );
  DFQD1 \mem_reg[71][8]  ( .D(n3525), .CP(clk), .Q(\mem[71][8] ) );
  DFQD1 \mem_reg[71][7]  ( .D(n3524), .CP(clk), .Q(\mem[71][7] ) );
  DFQD1 \mem_reg[71][6]  ( .D(n3523), .CP(clk), .Q(\mem[71][6] ) );
  DFQD1 \mem_reg[71][5]  ( .D(n3522), .CP(clk), .Q(\mem[71][5] ) );
  DFQD1 \mem_reg[71][4]  ( .D(n3521), .CP(clk), .Q(\mem[71][4] ) );
  DFQD1 \mem_reg[71][3]  ( .D(n3520), .CP(clk), .Q(\mem[71][3] ) );
  DFQD1 \mem_reg[71][2]  ( .D(n3519), .CP(clk), .Q(\mem[71][2] ) );
  DFQD1 \mem_reg[71][1]  ( .D(n3518), .CP(clk), .Q(\mem[71][1] ) );
  DFQD1 \mem_reg[71][0]  ( .D(n3517), .CP(clk), .Q(\mem[71][0] ) );
  DFQD1 \mem_reg[72][15]  ( .D(n3516), .CP(clk), .Q(\mem[72][15] ) );
  DFQD1 \mem_reg[72][14]  ( .D(n3515), .CP(clk), .Q(\mem[72][14] ) );
  DFQD1 \mem_reg[72][13]  ( .D(n3514), .CP(clk), .Q(\mem[72][13] ) );
  DFQD1 \mem_reg[72][12]  ( .D(n3513), .CP(clk), .Q(\mem[72][12] ) );
  DFQD1 \mem_reg[72][11]  ( .D(n3512), .CP(clk), .Q(\mem[72][11] ) );
  DFQD1 \mem_reg[72][10]  ( .D(n3511), .CP(clk), .Q(\mem[72][10] ) );
  DFQD1 \mem_reg[72][9]  ( .D(n3510), .CP(clk), .Q(\mem[72][9] ) );
  DFQD1 \mem_reg[72][8]  ( .D(n3509), .CP(clk), .Q(\mem[72][8] ) );
  DFQD1 \mem_reg[72][7]  ( .D(n3508), .CP(clk), .Q(\mem[72][7] ) );
  DFQD1 \mem_reg[72][6]  ( .D(n3507), .CP(clk), .Q(\mem[72][6] ) );
  DFQD1 \mem_reg[72][5]  ( .D(n3506), .CP(clk), .Q(\mem[72][5] ) );
  DFQD1 \mem_reg[72][4]  ( .D(n3505), .CP(clk), .Q(\mem[72][4] ) );
  DFQD1 \mem_reg[72][3]  ( .D(n3504), .CP(clk), .Q(\mem[72][3] ) );
  DFQD1 \mem_reg[72][2]  ( .D(n3503), .CP(clk), .Q(\mem[72][2] ) );
  DFQD1 \mem_reg[72][1]  ( .D(n3502), .CP(clk), .Q(\mem[72][1] ) );
  DFQD1 \mem_reg[72][0]  ( .D(n3501), .CP(clk), .Q(\mem[72][0] ) );
  DFQD1 \mem_reg[73][15]  ( .D(n3500), .CP(clk), .Q(\mem[73][15] ) );
  DFQD1 \mem_reg[73][14]  ( .D(n3499), .CP(clk), .Q(\mem[73][14] ) );
  DFQD1 \mem_reg[73][13]  ( .D(n3498), .CP(clk), .Q(\mem[73][13] ) );
  DFQD1 \mem_reg[73][12]  ( .D(n3497), .CP(clk), .Q(\mem[73][12] ) );
  DFQD1 \mem_reg[73][11]  ( .D(n3496), .CP(clk), .Q(\mem[73][11] ) );
  DFQD1 \mem_reg[73][10]  ( .D(n3495), .CP(clk), .Q(\mem[73][10] ) );
  DFQD1 \mem_reg[73][9]  ( .D(n3494), .CP(clk), .Q(\mem[73][9] ) );
  DFQD1 \mem_reg[73][8]  ( .D(n3493), .CP(clk), .Q(\mem[73][8] ) );
  DFQD1 \mem_reg[73][7]  ( .D(n3492), .CP(clk), .Q(\mem[73][7] ) );
  DFQD1 \mem_reg[73][6]  ( .D(n3491), .CP(clk), .Q(\mem[73][6] ) );
  DFQD1 \mem_reg[73][5]  ( .D(n3490), .CP(clk), .Q(\mem[73][5] ) );
  DFQD1 \mem_reg[73][4]  ( .D(n3489), .CP(clk), .Q(\mem[73][4] ) );
  DFQD1 \mem_reg[73][3]  ( .D(n3488), .CP(clk), .Q(\mem[73][3] ) );
  DFQD1 \mem_reg[73][2]  ( .D(n3487), .CP(clk), .Q(\mem[73][2] ) );
  DFQD1 \mem_reg[73][1]  ( .D(n3486), .CP(clk), .Q(\mem[73][1] ) );
  DFQD1 \mem_reg[73][0]  ( .D(n3485), .CP(clk), .Q(\mem[73][0] ) );
  DFQD1 \mem_reg[74][15]  ( .D(n3484), .CP(clk), .Q(\mem[74][15] ) );
  DFQD1 \mem_reg[74][14]  ( .D(n3483), .CP(clk), .Q(\mem[74][14] ) );
  DFQD1 \mem_reg[74][13]  ( .D(n3482), .CP(clk), .Q(\mem[74][13] ) );
  DFQD1 \mem_reg[74][12]  ( .D(n3481), .CP(clk), .Q(\mem[74][12] ) );
  DFQD1 \mem_reg[74][11]  ( .D(n3480), .CP(clk), .Q(\mem[74][11] ) );
  DFQD1 \mem_reg[74][10]  ( .D(n3479), .CP(clk), .Q(\mem[74][10] ) );
  DFQD1 \mem_reg[74][9]  ( .D(n3478), .CP(clk), .Q(\mem[74][9] ) );
  DFQD1 \mem_reg[74][8]  ( .D(n3477), .CP(clk), .Q(\mem[74][8] ) );
  DFQD1 \mem_reg[74][7]  ( .D(n3476), .CP(clk), .Q(\mem[74][7] ) );
  DFQD1 \mem_reg[74][6]  ( .D(n3475), .CP(clk), .Q(\mem[74][6] ) );
  DFQD1 \mem_reg[74][5]  ( .D(n3474), .CP(clk), .Q(\mem[74][5] ) );
  DFQD1 \mem_reg[74][4]  ( .D(n3473), .CP(clk), .Q(\mem[74][4] ) );
  DFQD1 \mem_reg[74][3]  ( .D(n3472), .CP(clk), .Q(\mem[74][3] ) );
  DFQD1 \mem_reg[74][2]  ( .D(n3471), .CP(clk), .Q(\mem[74][2] ) );
  DFQD1 \mem_reg[74][1]  ( .D(n3470), .CP(clk), .Q(\mem[74][1] ) );
  DFQD1 \mem_reg[74][0]  ( .D(n3469), .CP(clk), .Q(\mem[74][0] ) );
  DFQD1 \mem_reg[75][15]  ( .D(n3468), .CP(clk), .Q(\mem[75][15] ) );
  DFQD1 \mem_reg[75][14]  ( .D(n3467), .CP(clk), .Q(\mem[75][14] ) );
  DFQD1 \mem_reg[75][13]  ( .D(n3466), .CP(clk), .Q(\mem[75][13] ) );
  DFQD1 \mem_reg[75][12]  ( .D(n3465), .CP(clk), .Q(\mem[75][12] ) );
  DFQD1 \mem_reg[75][11]  ( .D(n3464), .CP(clk), .Q(\mem[75][11] ) );
  DFQD1 \mem_reg[75][10]  ( .D(n3463), .CP(clk), .Q(\mem[75][10] ) );
  DFQD1 \mem_reg[75][9]  ( .D(n3462), .CP(clk), .Q(\mem[75][9] ) );
  DFQD1 \mem_reg[75][8]  ( .D(n3461), .CP(clk), .Q(\mem[75][8] ) );
  DFQD1 \mem_reg[75][7]  ( .D(n3460), .CP(clk), .Q(\mem[75][7] ) );
  DFQD1 \mem_reg[75][6]  ( .D(n3459), .CP(clk), .Q(\mem[75][6] ) );
  DFQD1 \mem_reg[75][5]  ( .D(n3458), .CP(clk), .Q(\mem[75][5] ) );
  DFQD1 \mem_reg[75][4]  ( .D(n3457), .CP(clk), .Q(\mem[75][4] ) );
  DFQD1 \mem_reg[75][3]  ( .D(n3456), .CP(clk), .Q(\mem[75][3] ) );
  DFQD1 \mem_reg[75][2]  ( .D(n3455), .CP(clk), .Q(\mem[75][2] ) );
  DFQD1 \mem_reg[75][1]  ( .D(n3454), .CP(clk), .Q(\mem[75][1] ) );
  DFQD1 \mem_reg[75][0]  ( .D(n3453), .CP(clk), .Q(\mem[75][0] ) );
  DFQD1 \mem_reg[76][15]  ( .D(n3452), .CP(clk), .Q(\mem[76][15] ) );
  DFQD1 \mem_reg[76][14]  ( .D(n3451), .CP(clk), .Q(\mem[76][14] ) );
  DFQD1 \mem_reg[76][13]  ( .D(n3450), .CP(clk), .Q(\mem[76][13] ) );
  DFQD1 \mem_reg[76][12]  ( .D(n3449), .CP(clk), .Q(\mem[76][12] ) );
  DFQD1 \mem_reg[76][11]  ( .D(n3448), .CP(clk), .Q(\mem[76][11] ) );
  DFQD1 \mem_reg[76][10]  ( .D(n3447), .CP(clk), .Q(\mem[76][10] ) );
  DFQD1 \mem_reg[76][9]  ( .D(n3446), .CP(clk), .Q(\mem[76][9] ) );
  DFQD1 \mem_reg[76][8]  ( .D(n3445), .CP(clk), .Q(\mem[76][8] ) );
  DFQD1 \mem_reg[76][7]  ( .D(n3444), .CP(clk), .Q(\mem[76][7] ) );
  DFQD1 \mem_reg[76][6]  ( .D(n3443), .CP(clk), .Q(\mem[76][6] ) );
  DFQD1 \mem_reg[76][5]  ( .D(n3442), .CP(clk), .Q(\mem[76][5] ) );
  DFQD1 \mem_reg[76][4]  ( .D(n3441), .CP(clk), .Q(\mem[76][4] ) );
  DFQD1 \mem_reg[76][3]  ( .D(n3440), .CP(clk), .Q(\mem[76][3] ) );
  DFQD1 \mem_reg[76][2]  ( .D(n3439), .CP(clk), .Q(\mem[76][2] ) );
  DFQD1 \mem_reg[76][1]  ( .D(n3438), .CP(clk), .Q(\mem[76][1] ) );
  DFQD1 \mem_reg[76][0]  ( .D(n3437), .CP(clk), .Q(\mem[76][0] ) );
  DFQD1 \mem_reg[77][15]  ( .D(n3436), .CP(clk), .Q(\mem[77][15] ) );
  DFQD1 \mem_reg[77][14]  ( .D(n3435), .CP(clk), .Q(\mem[77][14] ) );
  DFQD1 \mem_reg[77][13]  ( .D(n3434), .CP(clk), .Q(\mem[77][13] ) );
  DFQD1 \mem_reg[77][12]  ( .D(n3433), .CP(clk), .Q(\mem[77][12] ) );
  DFQD1 \mem_reg[77][11]  ( .D(n3432), .CP(clk), .Q(\mem[77][11] ) );
  DFQD1 \mem_reg[77][10]  ( .D(n3431), .CP(clk), .Q(\mem[77][10] ) );
  DFQD1 \mem_reg[77][9]  ( .D(n3430), .CP(clk), .Q(\mem[77][9] ) );
  DFQD1 \mem_reg[77][8]  ( .D(n3429), .CP(clk), .Q(\mem[77][8] ) );
  DFQD1 \mem_reg[77][7]  ( .D(n3428), .CP(clk), .Q(\mem[77][7] ) );
  DFQD1 \mem_reg[77][6]  ( .D(n3427), .CP(clk), .Q(\mem[77][6] ) );
  DFQD1 \mem_reg[77][5]  ( .D(n3426), .CP(clk), .Q(\mem[77][5] ) );
  DFQD1 \mem_reg[77][4]  ( .D(n3425), .CP(clk), .Q(\mem[77][4] ) );
  DFQD1 \mem_reg[77][3]  ( .D(n3424), .CP(clk), .Q(\mem[77][3] ) );
  DFQD1 \mem_reg[77][2]  ( .D(n3423), .CP(clk), .Q(\mem[77][2] ) );
  DFQD1 \mem_reg[77][1]  ( .D(n3422), .CP(clk), .Q(\mem[77][1] ) );
  DFQD1 \mem_reg[77][0]  ( .D(n3421), .CP(clk), .Q(\mem[77][0] ) );
  DFQD1 \mem_reg[78][15]  ( .D(n3420), .CP(clk), .Q(\mem[78][15] ) );
  DFQD1 \mem_reg[78][14]  ( .D(n3419), .CP(clk), .Q(\mem[78][14] ) );
  DFQD1 \mem_reg[78][13]  ( .D(n3418), .CP(clk), .Q(\mem[78][13] ) );
  DFQD1 \mem_reg[78][12]  ( .D(n3417), .CP(clk), .Q(\mem[78][12] ) );
  DFQD1 \mem_reg[78][11]  ( .D(n3416), .CP(clk), .Q(\mem[78][11] ) );
  DFQD1 \mem_reg[78][10]  ( .D(n3415), .CP(clk), .Q(\mem[78][10] ) );
  DFQD1 \mem_reg[78][9]  ( .D(n3414), .CP(clk), .Q(\mem[78][9] ) );
  DFQD1 \mem_reg[78][8]  ( .D(n3413), .CP(clk), .Q(\mem[78][8] ) );
  DFQD1 \mem_reg[78][7]  ( .D(n3412), .CP(clk), .Q(\mem[78][7] ) );
  DFQD1 \mem_reg[78][6]  ( .D(n3411), .CP(clk), .Q(\mem[78][6] ) );
  DFQD1 \mem_reg[78][5]  ( .D(n3410), .CP(clk), .Q(\mem[78][5] ) );
  DFQD1 \mem_reg[78][4]  ( .D(n3409), .CP(clk), .Q(\mem[78][4] ) );
  DFQD1 \mem_reg[78][3]  ( .D(n3408), .CP(clk), .Q(\mem[78][3] ) );
  DFQD1 \mem_reg[78][2]  ( .D(n3407), .CP(clk), .Q(\mem[78][2] ) );
  DFQD1 \mem_reg[78][1]  ( .D(n3406), .CP(clk), .Q(\mem[78][1] ) );
  DFQD1 \mem_reg[78][0]  ( .D(n3405), .CP(clk), .Q(\mem[78][0] ) );
  DFQD1 \mem_reg[79][15]  ( .D(n3404), .CP(clk), .Q(\mem[79][15] ) );
  DFQD1 \mem_reg[79][14]  ( .D(n3403), .CP(clk), .Q(\mem[79][14] ) );
  DFQD1 \mem_reg[79][13]  ( .D(n3402), .CP(clk), .Q(\mem[79][13] ) );
  DFQD1 \mem_reg[79][12]  ( .D(n3401), .CP(clk), .Q(\mem[79][12] ) );
  DFQD1 \mem_reg[79][11]  ( .D(n3400), .CP(clk), .Q(\mem[79][11] ) );
  DFQD1 \mem_reg[79][10]  ( .D(n3399), .CP(clk), .Q(\mem[79][10] ) );
  DFQD1 \mem_reg[79][9]  ( .D(n3398), .CP(clk), .Q(\mem[79][9] ) );
  DFQD1 \mem_reg[79][8]  ( .D(n3397), .CP(clk), .Q(\mem[79][8] ) );
  DFQD1 \mem_reg[79][7]  ( .D(n3396), .CP(clk), .Q(\mem[79][7] ) );
  DFQD1 \mem_reg[79][6]  ( .D(n3395), .CP(clk), .Q(\mem[79][6] ) );
  DFQD1 \mem_reg[79][5]  ( .D(n3394), .CP(clk), .Q(\mem[79][5] ) );
  DFQD1 \mem_reg[79][4]  ( .D(n3393), .CP(clk), .Q(\mem[79][4] ) );
  DFQD1 \mem_reg[79][3]  ( .D(n3392), .CP(clk), .Q(\mem[79][3] ) );
  DFQD1 \mem_reg[79][2]  ( .D(n3391), .CP(clk), .Q(\mem[79][2] ) );
  DFQD1 \mem_reg[79][1]  ( .D(n3390), .CP(clk), .Q(\mem[79][1] ) );
  DFQD1 \mem_reg[79][0]  ( .D(n3389), .CP(clk), .Q(\mem[79][0] ) );
  DFQD1 \mem_reg[80][15]  ( .D(n3388), .CP(clk), .Q(\mem[80][15] ) );
  DFQD1 \mem_reg[80][14]  ( .D(n3387), .CP(clk), .Q(\mem[80][14] ) );
  DFQD1 \mem_reg[80][13]  ( .D(n3386), .CP(clk), .Q(\mem[80][13] ) );
  DFQD1 \mem_reg[80][12]  ( .D(n3385), .CP(clk), .Q(\mem[80][12] ) );
  DFQD1 \mem_reg[80][11]  ( .D(n3384), .CP(clk), .Q(\mem[80][11] ) );
  DFQD1 \mem_reg[80][10]  ( .D(n3383), .CP(clk), .Q(\mem[80][10] ) );
  DFQD1 \mem_reg[80][9]  ( .D(n3382), .CP(clk), .Q(\mem[80][9] ) );
  DFQD1 \mem_reg[80][8]  ( .D(n3381), .CP(clk), .Q(\mem[80][8] ) );
  DFQD1 \mem_reg[80][7]  ( .D(n3380), .CP(clk), .Q(\mem[80][7] ) );
  DFQD1 \mem_reg[80][6]  ( .D(n3379), .CP(clk), .Q(\mem[80][6] ) );
  DFQD1 \mem_reg[80][5]  ( .D(n3378), .CP(clk), .Q(\mem[80][5] ) );
  DFQD1 \mem_reg[80][4]  ( .D(n3377), .CP(clk), .Q(\mem[80][4] ) );
  DFQD1 \mem_reg[80][3]  ( .D(n3376), .CP(clk), .Q(\mem[80][3] ) );
  DFQD1 \mem_reg[80][2]  ( .D(n3375), .CP(clk), .Q(\mem[80][2] ) );
  DFQD1 \mem_reg[80][1]  ( .D(n3374), .CP(clk), .Q(\mem[80][1] ) );
  DFQD1 \mem_reg[80][0]  ( .D(n3373), .CP(clk), .Q(\mem[80][0] ) );
  DFQD1 \mem_reg[81][15]  ( .D(n3372), .CP(clk), .Q(\mem[81][15] ) );
  DFQD1 \mem_reg[81][14]  ( .D(n3371), .CP(clk), .Q(\mem[81][14] ) );
  DFQD1 \mem_reg[81][13]  ( .D(n3370), .CP(clk), .Q(\mem[81][13] ) );
  DFQD1 \mem_reg[81][12]  ( .D(n3369), .CP(clk), .Q(\mem[81][12] ) );
  DFQD1 \mem_reg[81][11]  ( .D(n3368), .CP(clk), .Q(\mem[81][11] ) );
  DFQD1 \mem_reg[81][10]  ( .D(n3367), .CP(clk), .Q(\mem[81][10] ) );
  DFQD1 \mem_reg[81][9]  ( .D(n3366), .CP(clk), .Q(\mem[81][9] ) );
  DFQD1 \mem_reg[81][8]  ( .D(n3365), .CP(clk), .Q(\mem[81][8] ) );
  DFQD1 \mem_reg[81][7]  ( .D(n3364), .CP(clk), .Q(\mem[81][7] ) );
  DFQD1 \mem_reg[81][6]  ( .D(n3363), .CP(clk), .Q(\mem[81][6] ) );
  DFQD1 \mem_reg[81][5]  ( .D(n3362), .CP(clk), .Q(\mem[81][5] ) );
  DFQD1 \mem_reg[81][4]  ( .D(n3361), .CP(clk), .Q(\mem[81][4] ) );
  DFQD1 \mem_reg[81][3]  ( .D(n3360), .CP(clk), .Q(\mem[81][3] ) );
  DFQD1 \mem_reg[81][2]  ( .D(n3359), .CP(clk), .Q(\mem[81][2] ) );
  DFQD1 \mem_reg[81][1]  ( .D(n3358), .CP(clk), .Q(\mem[81][1] ) );
  DFQD1 \mem_reg[81][0]  ( .D(n3357), .CP(clk), .Q(\mem[81][0] ) );
  DFQD1 \mem_reg[82][15]  ( .D(n3356), .CP(clk), .Q(\mem[82][15] ) );
  DFQD1 \mem_reg[82][14]  ( .D(n3355), .CP(clk), .Q(\mem[82][14] ) );
  DFQD1 \mem_reg[82][13]  ( .D(n3354), .CP(clk), .Q(\mem[82][13] ) );
  DFQD1 \mem_reg[82][12]  ( .D(n3353), .CP(clk), .Q(\mem[82][12] ) );
  DFQD1 \mem_reg[82][11]  ( .D(n3352), .CP(clk), .Q(\mem[82][11] ) );
  DFQD1 \mem_reg[82][10]  ( .D(n3351), .CP(clk), .Q(\mem[82][10] ) );
  DFQD1 \mem_reg[82][9]  ( .D(n3350), .CP(clk), .Q(\mem[82][9] ) );
  DFQD1 \mem_reg[82][8]  ( .D(n3349), .CP(clk), .Q(\mem[82][8] ) );
  DFQD1 \mem_reg[82][7]  ( .D(n3348), .CP(clk), .Q(\mem[82][7] ) );
  DFQD1 \mem_reg[82][6]  ( .D(n3347), .CP(clk), .Q(\mem[82][6] ) );
  DFQD1 \mem_reg[82][5]  ( .D(n3346), .CP(clk), .Q(\mem[82][5] ) );
  DFQD1 \mem_reg[82][4]  ( .D(n3345), .CP(clk), .Q(\mem[82][4] ) );
  DFQD1 \mem_reg[82][3]  ( .D(n3344), .CP(clk), .Q(\mem[82][3] ) );
  DFQD1 \mem_reg[82][2]  ( .D(n3343), .CP(clk), .Q(\mem[82][2] ) );
  DFQD1 \mem_reg[82][1]  ( .D(n3342), .CP(clk), .Q(\mem[82][1] ) );
  DFQD1 \mem_reg[82][0]  ( .D(n3341), .CP(clk), .Q(\mem[82][0] ) );
  DFQD1 \mem_reg[83][15]  ( .D(n3340), .CP(clk), .Q(\mem[83][15] ) );
  DFQD1 \mem_reg[83][14]  ( .D(n3339), .CP(clk), .Q(\mem[83][14] ) );
  DFQD1 \mem_reg[83][13]  ( .D(n3338), .CP(clk), .Q(\mem[83][13] ) );
  DFQD1 \mem_reg[83][12]  ( .D(n3337), .CP(clk), .Q(\mem[83][12] ) );
  DFQD1 \mem_reg[83][11]  ( .D(n3336), .CP(clk), .Q(\mem[83][11] ) );
  DFQD1 \mem_reg[83][10]  ( .D(n3335), .CP(clk), .Q(\mem[83][10] ) );
  DFQD1 \mem_reg[83][9]  ( .D(n3334), .CP(clk), .Q(\mem[83][9] ) );
  DFQD1 \mem_reg[83][8]  ( .D(n3333), .CP(clk), .Q(\mem[83][8] ) );
  DFQD1 \mem_reg[83][7]  ( .D(n3332), .CP(clk), .Q(\mem[83][7] ) );
  DFQD1 \mem_reg[83][6]  ( .D(n3331), .CP(clk), .Q(\mem[83][6] ) );
  DFQD1 \mem_reg[83][5]  ( .D(n3330), .CP(clk), .Q(\mem[83][5] ) );
  DFQD1 \mem_reg[83][4]  ( .D(n3329), .CP(clk), .Q(\mem[83][4] ) );
  DFQD1 \mem_reg[83][3]  ( .D(n3328), .CP(clk), .Q(\mem[83][3] ) );
  DFQD1 \mem_reg[83][2]  ( .D(n3327), .CP(clk), .Q(\mem[83][2] ) );
  DFQD1 \mem_reg[83][1]  ( .D(n3326), .CP(clk), .Q(\mem[83][1] ) );
  DFQD1 \mem_reg[83][0]  ( .D(n3325), .CP(clk), .Q(\mem[83][0] ) );
  DFQD1 \mem_reg[84][15]  ( .D(n3324), .CP(clk), .Q(\mem[84][15] ) );
  DFQD1 \mem_reg[84][14]  ( .D(n3323), .CP(clk), .Q(\mem[84][14] ) );
  DFQD1 \mem_reg[84][13]  ( .D(n3322), .CP(clk), .Q(\mem[84][13] ) );
  DFQD1 \mem_reg[84][12]  ( .D(n3321), .CP(clk), .Q(\mem[84][12] ) );
  DFQD1 \mem_reg[84][11]  ( .D(n3320), .CP(clk), .Q(\mem[84][11] ) );
  DFQD1 \mem_reg[84][10]  ( .D(n3319), .CP(clk), .Q(\mem[84][10] ) );
  DFQD1 \mem_reg[84][9]  ( .D(n3318), .CP(clk), .Q(\mem[84][9] ) );
  DFQD1 \mem_reg[84][8]  ( .D(n3317), .CP(clk), .Q(\mem[84][8] ) );
  DFQD1 \mem_reg[84][7]  ( .D(n3316), .CP(clk), .Q(\mem[84][7] ) );
  DFQD1 \mem_reg[84][6]  ( .D(n3315), .CP(clk), .Q(\mem[84][6] ) );
  DFQD1 \mem_reg[84][5]  ( .D(n3314), .CP(clk), .Q(\mem[84][5] ) );
  DFQD1 \mem_reg[84][4]  ( .D(n3313), .CP(clk), .Q(\mem[84][4] ) );
  DFQD1 \mem_reg[84][3]  ( .D(n3312), .CP(clk), .Q(\mem[84][3] ) );
  DFQD1 \mem_reg[84][2]  ( .D(n3311), .CP(clk), .Q(\mem[84][2] ) );
  DFQD1 \mem_reg[84][1]  ( .D(n3310), .CP(clk), .Q(\mem[84][1] ) );
  DFQD1 \mem_reg[84][0]  ( .D(n3309), .CP(clk), .Q(\mem[84][0] ) );
  DFQD1 \mem_reg[85][15]  ( .D(n3308), .CP(clk), .Q(\mem[85][15] ) );
  DFQD1 \mem_reg[85][14]  ( .D(n3307), .CP(clk), .Q(\mem[85][14] ) );
  DFQD1 \mem_reg[85][13]  ( .D(n3306), .CP(clk), .Q(\mem[85][13] ) );
  DFQD1 \mem_reg[85][12]  ( .D(n3305), .CP(clk), .Q(\mem[85][12] ) );
  DFQD1 \mem_reg[85][11]  ( .D(n3304), .CP(clk), .Q(\mem[85][11] ) );
  DFQD1 \mem_reg[85][10]  ( .D(n3303), .CP(clk), .Q(\mem[85][10] ) );
  DFQD1 \mem_reg[85][9]  ( .D(n3302), .CP(clk), .Q(\mem[85][9] ) );
  DFQD1 \mem_reg[85][8]  ( .D(n3301), .CP(clk), .Q(\mem[85][8] ) );
  DFQD1 \mem_reg[85][7]  ( .D(n3300), .CP(clk), .Q(\mem[85][7] ) );
  DFQD1 \mem_reg[85][6]  ( .D(n3299), .CP(clk), .Q(\mem[85][6] ) );
  DFQD1 \mem_reg[85][5]  ( .D(n3298), .CP(clk), .Q(\mem[85][5] ) );
  DFQD1 \mem_reg[85][4]  ( .D(n3297), .CP(clk), .Q(\mem[85][4] ) );
  DFQD1 \mem_reg[85][3]  ( .D(n3296), .CP(clk), .Q(\mem[85][3] ) );
  DFQD1 \mem_reg[85][2]  ( .D(n3295), .CP(clk), .Q(\mem[85][2] ) );
  DFQD1 \mem_reg[85][1]  ( .D(n3294), .CP(clk), .Q(\mem[85][1] ) );
  DFQD1 \mem_reg[85][0]  ( .D(n3293), .CP(clk), .Q(\mem[85][0] ) );
  DFQD1 \mem_reg[86][15]  ( .D(n3292), .CP(clk), .Q(\mem[86][15] ) );
  DFQD1 \mem_reg[86][14]  ( .D(n3291), .CP(clk), .Q(\mem[86][14] ) );
  DFQD1 \mem_reg[86][13]  ( .D(n3290), .CP(clk), .Q(\mem[86][13] ) );
  DFQD1 \mem_reg[86][12]  ( .D(n3289), .CP(clk), .Q(\mem[86][12] ) );
  DFQD1 \mem_reg[86][11]  ( .D(n3288), .CP(clk), .Q(\mem[86][11] ) );
  DFQD1 \mem_reg[86][10]  ( .D(n3287), .CP(clk), .Q(\mem[86][10] ) );
  DFQD1 \mem_reg[86][9]  ( .D(n3286), .CP(clk), .Q(\mem[86][9] ) );
  DFQD1 \mem_reg[86][8]  ( .D(n3285), .CP(clk), .Q(\mem[86][8] ) );
  DFQD1 \mem_reg[86][7]  ( .D(n3284), .CP(clk), .Q(\mem[86][7] ) );
  DFQD1 \mem_reg[86][6]  ( .D(n3283), .CP(clk), .Q(\mem[86][6] ) );
  DFQD1 \mem_reg[86][5]  ( .D(n3282), .CP(clk), .Q(\mem[86][5] ) );
  DFQD1 \mem_reg[86][4]  ( .D(n3281), .CP(clk), .Q(\mem[86][4] ) );
  DFQD1 \mem_reg[86][3]  ( .D(n3280), .CP(clk), .Q(\mem[86][3] ) );
  DFQD1 \mem_reg[86][2]  ( .D(n3279), .CP(clk), .Q(\mem[86][2] ) );
  DFQD1 \mem_reg[86][1]  ( .D(n3278), .CP(clk), .Q(\mem[86][1] ) );
  DFQD1 \mem_reg[86][0]  ( .D(n3277), .CP(clk), .Q(\mem[86][0] ) );
  DFQD1 \mem_reg[87][15]  ( .D(n3276), .CP(clk), .Q(\mem[87][15] ) );
  DFQD1 \mem_reg[87][14]  ( .D(n3275), .CP(clk), .Q(\mem[87][14] ) );
  DFQD1 \mem_reg[87][13]  ( .D(n3274), .CP(clk), .Q(\mem[87][13] ) );
  DFQD1 \mem_reg[87][12]  ( .D(n3273), .CP(clk), .Q(\mem[87][12] ) );
  DFQD1 \mem_reg[87][11]  ( .D(n3272), .CP(clk), .Q(\mem[87][11] ) );
  DFQD1 \mem_reg[87][10]  ( .D(n3271), .CP(clk), .Q(\mem[87][10] ) );
  DFQD1 \mem_reg[87][9]  ( .D(n3270), .CP(clk), .Q(\mem[87][9] ) );
  DFQD1 \mem_reg[87][8]  ( .D(n3269), .CP(clk), .Q(\mem[87][8] ) );
  DFQD1 \mem_reg[87][7]  ( .D(n3268), .CP(clk), .Q(\mem[87][7] ) );
  DFQD1 \mem_reg[87][6]  ( .D(n3267), .CP(clk), .Q(\mem[87][6] ) );
  DFQD1 \mem_reg[87][5]  ( .D(n3266), .CP(clk), .Q(\mem[87][5] ) );
  DFQD1 \mem_reg[87][4]  ( .D(n3265), .CP(clk), .Q(\mem[87][4] ) );
  DFQD1 \mem_reg[87][3]  ( .D(n3264), .CP(clk), .Q(\mem[87][3] ) );
  DFQD1 \mem_reg[87][2]  ( .D(n3263), .CP(clk), .Q(\mem[87][2] ) );
  DFQD1 \mem_reg[87][1]  ( .D(n3262), .CP(clk), .Q(\mem[87][1] ) );
  DFQD1 \mem_reg[87][0]  ( .D(n3261), .CP(clk), .Q(\mem[87][0] ) );
  DFQD1 \mem_reg[88][15]  ( .D(n3260), .CP(clk), .Q(\mem[88][15] ) );
  DFQD1 \mem_reg[88][14]  ( .D(n3259), .CP(clk), .Q(\mem[88][14] ) );
  DFQD1 \mem_reg[88][13]  ( .D(n3258), .CP(clk), .Q(\mem[88][13] ) );
  DFQD1 \mem_reg[88][12]  ( .D(n3257), .CP(clk), .Q(\mem[88][12] ) );
  DFQD1 \mem_reg[88][11]  ( .D(n3256), .CP(clk), .Q(\mem[88][11] ) );
  DFQD1 \mem_reg[88][10]  ( .D(n3255), .CP(clk), .Q(\mem[88][10] ) );
  DFQD1 \mem_reg[88][9]  ( .D(n3254), .CP(clk), .Q(\mem[88][9] ) );
  DFQD1 \mem_reg[88][8]  ( .D(n3253), .CP(clk), .Q(\mem[88][8] ) );
  DFQD1 \mem_reg[88][7]  ( .D(n3252), .CP(clk), .Q(\mem[88][7] ) );
  DFQD1 \mem_reg[88][6]  ( .D(n3251), .CP(clk), .Q(\mem[88][6] ) );
  DFQD1 \mem_reg[88][5]  ( .D(n3250), .CP(clk), .Q(\mem[88][5] ) );
  DFQD1 \mem_reg[88][4]  ( .D(n3249), .CP(clk), .Q(\mem[88][4] ) );
  DFQD1 \mem_reg[88][3]  ( .D(n3248), .CP(clk), .Q(\mem[88][3] ) );
  DFQD1 \mem_reg[88][2]  ( .D(n3247), .CP(clk), .Q(\mem[88][2] ) );
  DFQD1 \mem_reg[88][1]  ( .D(n3246), .CP(clk), .Q(\mem[88][1] ) );
  DFQD1 \mem_reg[88][0]  ( .D(n3245), .CP(clk), .Q(\mem[88][0] ) );
  DFQD1 \mem_reg[89][15]  ( .D(n3244), .CP(clk), .Q(\mem[89][15] ) );
  DFQD1 \mem_reg[89][14]  ( .D(n3243), .CP(clk), .Q(\mem[89][14] ) );
  DFQD1 \mem_reg[89][13]  ( .D(n3242), .CP(clk), .Q(\mem[89][13] ) );
  DFQD1 \mem_reg[89][12]  ( .D(n3241), .CP(clk), .Q(\mem[89][12] ) );
  DFQD1 \mem_reg[89][11]  ( .D(n3240), .CP(clk), .Q(\mem[89][11] ) );
  DFQD1 \mem_reg[89][10]  ( .D(n3239), .CP(clk), .Q(\mem[89][10] ) );
  DFQD1 \mem_reg[89][9]  ( .D(n3238), .CP(clk), .Q(\mem[89][9] ) );
  DFQD1 \mem_reg[89][8]  ( .D(n3237), .CP(clk), .Q(\mem[89][8] ) );
  DFQD1 \mem_reg[89][7]  ( .D(n3236), .CP(clk), .Q(\mem[89][7] ) );
  DFQD1 \mem_reg[89][6]  ( .D(n3235), .CP(clk), .Q(\mem[89][6] ) );
  DFQD1 \mem_reg[89][5]  ( .D(n3234), .CP(clk), .Q(\mem[89][5] ) );
  DFQD1 \mem_reg[89][4]  ( .D(n3233), .CP(clk), .Q(\mem[89][4] ) );
  DFQD1 \mem_reg[89][3]  ( .D(n3232), .CP(clk), .Q(\mem[89][3] ) );
  DFQD1 \mem_reg[89][2]  ( .D(n3231), .CP(clk), .Q(\mem[89][2] ) );
  DFQD1 \mem_reg[89][1]  ( .D(n3230), .CP(clk), .Q(\mem[89][1] ) );
  DFQD1 \mem_reg[89][0]  ( .D(n3229), .CP(clk), .Q(\mem[89][0] ) );
  DFQD1 \mem_reg[90][15]  ( .D(n3228), .CP(clk), .Q(\mem[90][15] ) );
  DFQD1 \mem_reg[90][14]  ( .D(n3227), .CP(clk), .Q(\mem[90][14] ) );
  DFQD1 \mem_reg[90][13]  ( .D(n3226), .CP(clk), .Q(\mem[90][13] ) );
  DFQD1 \mem_reg[90][12]  ( .D(n3225), .CP(clk), .Q(\mem[90][12] ) );
  DFQD1 \mem_reg[90][11]  ( .D(n3224), .CP(clk), .Q(\mem[90][11] ) );
  DFQD1 \mem_reg[90][10]  ( .D(n3223), .CP(clk), .Q(\mem[90][10] ) );
  DFQD1 \mem_reg[90][9]  ( .D(n3222), .CP(clk), .Q(\mem[90][9] ) );
  DFQD1 \mem_reg[90][8]  ( .D(n3221), .CP(clk), .Q(\mem[90][8] ) );
  DFQD1 \mem_reg[90][7]  ( .D(n3220), .CP(clk), .Q(\mem[90][7] ) );
  DFQD1 \mem_reg[90][6]  ( .D(n3219), .CP(clk), .Q(\mem[90][6] ) );
  DFQD1 \mem_reg[90][5]  ( .D(n3218), .CP(clk), .Q(\mem[90][5] ) );
  DFQD1 \mem_reg[90][4]  ( .D(n3217), .CP(clk), .Q(\mem[90][4] ) );
  DFQD1 \mem_reg[90][3]  ( .D(n3216), .CP(clk), .Q(\mem[90][3] ) );
  DFQD1 \mem_reg[90][2]  ( .D(n3215), .CP(clk), .Q(\mem[90][2] ) );
  DFQD1 \mem_reg[90][1]  ( .D(n3214), .CP(clk), .Q(\mem[90][1] ) );
  DFQD1 \mem_reg[90][0]  ( .D(n3213), .CP(clk), .Q(\mem[90][0] ) );
  DFQD1 \mem_reg[91][15]  ( .D(n3212), .CP(clk), .Q(\mem[91][15] ) );
  DFQD1 \mem_reg[91][14]  ( .D(n3211), .CP(clk), .Q(\mem[91][14] ) );
  DFQD1 \mem_reg[91][13]  ( .D(n3210), .CP(clk), .Q(\mem[91][13] ) );
  DFQD1 \mem_reg[91][12]  ( .D(n3209), .CP(clk), .Q(\mem[91][12] ) );
  DFQD1 \mem_reg[91][11]  ( .D(n3208), .CP(clk), .Q(\mem[91][11] ) );
  DFQD1 \mem_reg[91][10]  ( .D(n3207), .CP(clk), .Q(\mem[91][10] ) );
  DFQD1 \mem_reg[91][9]  ( .D(n3206), .CP(clk), .Q(\mem[91][9] ) );
  DFQD1 \mem_reg[91][8]  ( .D(n3205), .CP(clk), .Q(\mem[91][8] ) );
  DFQD1 \mem_reg[91][7]  ( .D(n3204), .CP(clk), .Q(\mem[91][7] ) );
  DFQD1 \mem_reg[91][6]  ( .D(n3203), .CP(clk), .Q(\mem[91][6] ) );
  DFQD1 \mem_reg[91][5]  ( .D(n3202), .CP(clk), .Q(\mem[91][5] ) );
  DFQD1 \mem_reg[91][4]  ( .D(n3201), .CP(clk), .Q(\mem[91][4] ) );
  DFQD1 \mem_reg[91][3]  ( .D(n3200), .CP(clk), .Q(\mem[91][3] ) );
  DFQD1 \mem_reg[91][2]  ( .D(n3199), .CP(clk), .Q(\mem[91][2] ) );
  DFQD1 \mem_reg[91][1]  ( .D(n3198), .CP(clk), .Q(\mem[91][1] ) );
  DFQD1 \mem_reg[91][0]  ( .D(n3197), .CP(clk), .Q(\mem[91][0] ) );
  DFQD1 \mem_reg[92][15]  ( .D(n3196), .CP(clk), .Q(\mem[92][15] ) );
  DFQD1 \mem_reg[92][14]  ( .D(n3195), .CP(clk), .Q(\mem[92][14] ) );
  DFQD1 \mem_reg[92][13]  ( .D(n3194), .CP(clk), .Q(\mem[92][13] ) );
  DFQD1 \mem_reg[92][12]  ( .D(n3193), .CP(clk), .Q(\mem[92][12] ) );
  DFQD1 \mem_reg[92][11]  ( .D(n3192), .CP(clk), .Q(\mem[92][11] ) );
  DFQD1 \mem_reg[92][10]  ( .D(n3191), .CP(clk), .Q(\mem[92][10] ) );
  DFQD1 \mem_reg[92][9]  ( .D(n3190), .CP(clk), .Q(\mem[92][9] ) );
  DFQD1 \mem_reg[92][8]  ( .D(n3189), .CP(clk), .Q(\mem[92][8] ) );
  DFQD1 \mem_reg[92][7]  ( .D(n3188), .CP(clk), .Q(\mem[92][7] ) );
  DFQD1 \mem_reg[92][6]  ( .D(n3187), .CP(clk), .Q(\mem[92][6] ) );
  DFQD1 \mem_reg[92][5]  ( .D(n3186), .CP(clk), .Q(\mem[92][5] ) );
  DFQD1 \mem_reg[92][4]  ( .D(n3185), .CP(clk), .Q(\mem[92][4] ) );
  DFQD1 \mem_reg[92][3]  ( .D(n3184), .CP(clk), .Q(\mem[92][3] ) );
  DFQD1 \mem_reg[92][2]  ( .D(n3183), .CP(clk), .Q(\mem[92][2] ) );
  DFQD1 \mem_reg[92][1]  ( .D(n3182), .CP(clk), .Q(\mem[92][1] ) );
  DFQD1 \mem_reg[92][0]  ( .D(n3181), .CP(clk), .Q(\mem[92][0] ) );
  DFQD1 \mem_reg[93][15]  ( .D(n3180), .CP(clk), .Q(\mem[93][15] ) );
  DFQD1 \mem_reg[93][14]  ( .D(n3179), .CP(clk), .Q(\mem[93][14] ) );
  DFQD1 \mem_reg[93][13]  ( .D(n3178), .CP(clk), .Q(\mem[93][13] ) );
  DFQD1 \mem_reg[93][12]  ( .D(n3177), .CP(clk), .Q(\mem[93][12] ) );
  DFQD1 \mem_reg[93][11]  ( .D(n3176), .CP(clk), .Q(\mem[93][11] ) );
  DFQD1 \mem_reg[93][10]  ( .D(n3175), .CP(clk), .Q(\mem[93][10] ) );
  DFQD1 \mem_reg[93][9]  ( .D(n3174), .CP(clk), .Q(\mem[93][9] ) );
  DFQD1 \mem_reg[93][8]  ( .D(n3173), .CP(clk), .Q(\mem[93][8] ) );
  DFQD1 \mem_reg[93][7]  ( .D(n3172), .CP(clk), .Q(\mem[93][7] ) );
  DFQD1 \mem_reg[93][6]  ( .D(n3171), .CP(clk), .Q(\mem[93][6] ) );
  DFQD1 \mem_reg[93][5]  ( .D(n3170), .CP(clk), .Q(\mem[93][5] ) );
  DFQD1 \mem_reg[93][4]  ( .D(n3169), .CP(clk), .Q(\mem[93][4] ) );
  DFQD1 \mem_reg[93][3]  ( .D(n3168), .CP(clk), .Q(\mem[93][3] ) );
  DFQD1 \mem_reg[93][2]  ( .D(n3167), .CP(clk), .Q(\mem[93][2] ) );
  DFQD1 \mem_reg[93][1]  ( .D(n3166), .CP(clk), .Q(\mem[93][1] ) );
  DFQD1 \mem_reg[93][0]  ( .D(n3165), .CP(clk), .Q(\mem[93][0] ) );
  DFQD1 \mem_reg[94][15]  ( .D(n3164), .CP(clk), .Q(\mem[94][15] ) );
  DFQD1 \mem_reg[94][14]  ( .D(n3163), .CP(clk), .Q(\mem[94][14] ) );
  DFQD1 \mem_reg[94][13]  ( .D(n3162), .CP(clk), .Q(\mem[94][13] ) );
  DFQD1 \mem_reg[94][12]  ( .D(n3161), .CP(clk), .Q(\mem[94][12] ) );
  DFQD1 \mem_reg[94][11]  ( .D(n3160), .CP(clk), .Q(\mem[94][11] ) );
  DFQD1 \mem_reg[94][10]  ( .D(n3159), .CP(clk), .Q(\mem[94][10] ) );
  DFQD1 \mem_reg[94][9]  ( .D(n3158), .CP(clk), .Q(\mem[94][9] ) );
  DFQD1 \mem_reg[94][8]  ( .D(n3157), .CP(clk), .Q(\mem[94][8] ) );
  DFQD1 \mem_reg[94][7]  ( .D(n3156), .CP(clk), .Q(\mem[94][7] ) );
  DFQD1 \mem_reg[94][6]  ( .D(n3155), .CP(clk), .Q(\mem[94][6] ) );
  DFQD1 \mem_reg[94][5]  ( .D(n3154), .CP(clk), .Q(\mem[94][5] ) );
  DFQD1 \mem_reg[94][4]  ( .D(n3153), .CP(clk), .Q(\mem[94][4] ) );
  DFQD1 \mem_reg[94][3]  ( .D(n3152), .CP(clk), .Q(\mem[94][3] ) );
  DFQD1 \mem_reg[94][2]  ( .D(n3151), .CP(clk), .Q(\mem[94][2] ) );
  DFQD1 \mem_reg[94][1]  ( .D(n3150), .CP(clk), .Q(\mem[94][1] ) );
  DFQD1 \mem_reg[94][0]  ( .D(n3149), .CP(clk), .Q(\mem[94][0] ) );
  DFQD1 \mem_reg[95][15]  ( .D(n3148), .CP(clk), .Q(\mem[95][15] ) );
  DFQD1 \mem_reg[95][14]  ( .D(n3147), .CP(clk), .Q(\mem[95][14] ) );
  DFQD1 \mem_reg[95][13]  ( .D(n3146), .CP(clk), .Q(\mem[95][13] ) );
  DFQD1 \mem_reg[95][12]  ( .D(n3145), .CP(clk), .Q(\mem[95][12] ) );
  DFQD1 \mem_reg[95][11]  ( .D(n3144), .CP(clk), .Q(\mem[95][11] ) );
  DFQD1 \mem_reg[95][10]  ( .D(n3143), .CP(clk), .Q(\mem[95][10] ) );
  DFQD1 \mem_reg[95][9]  ( .D(n3142), .CP(clk), .Q(\mem[95][9] ) );
  DFQD1 \mem_reg[95][8]  ( .D(n3141), .CP(clk), .Q(\mem[95][8] ) );
  DFQD1 \mem_reg[95][7]  ( .D(n3140), .CP(clk), .Q(\mem[95][7] ) );
  DFQD1 \mem_reg[95][6]  ( .D(n3139), .CP(clk), .Q(\mem[95][6] ) );
  DFQD1 \mem_reg[95][5]  ( .D(n3138), .CP(clk), .Q(\mem[95][5] ) );
  DFQD1 \mem_reg[95][4]  ( .D(n3137), .CP(clk), .Q(\mem[95][4] ) );
  DFQD1 \mem_reg[95][3]  ( .D(n3136), .CP(clk), .Q(\mem[95][3] ) );
  DFQD1 \mem_reg[95][2]  ( .D(n3135), .CP(clk), .Q(\mem[95][2] ) );
  DFQD1 \mem_reg[95][1]  ( .D(n3134), .CP(clk), .Q(\mem[95][1] ) );
  DFQD1 \mem_reg[95][0]  ( .D(n3133), .CP(clk), .Q(\mem[95][0] ) );
  DFQD1 \mem_reg[96][15]  ( .D(n3132), .CP(clk), .Q(\mem[96][15] ) );
  DFQD1 \mem_reg[96][14]  ( .D(n3131), .CP(clk), .Q(\mem[96][14] ) );
  DFQD1 \mem_reg[96][13]  ( .D(n3130), .CP(clk), .Q(\mem[96][13] ) );
  DFQD1 \mem_reg[96][12]  ( .D(n3129), .CP(clk), .Q(\mem[96][12] ) );
  DFQD1 \mem_reg[96][11]  ( .D(n3128), .CP(clk), .Q(\mem[96][11] ) );
  DFQD1 \mem_reg[96][10]  ( .D(n3127), .CP(clk), .Q(\mem[96][10] ) );
  DFQD1 \mem_reg[96][9]  ( .D(n3126), .CP(clk), .Q(\mem[96][9] ) );
  DFQD1 \mem_reg[96][8]  ( .D(n3125), .CP(clk), .Q(\mem[96][8] ) );
  DFQD1 \mem_reg[96][7]  ( .D(n3124), .CP(clk), .Q(\mem[96][7] ) );
  DFQD1 \mem_reg[96][6]  ( .D(n3123), .CP(clk), .Q(\mem[96][6] ) );
  DFQD1 \mem_reg[96][5]  ( .D(n3122), .CP(clk), .Q(\mem[96][5] ) );
  DFQD1 \mem_reg[96][4]  ( .D(n3121), .CP(clk), .Q(\mem[96][4] ) );
  DFQD1 \mem_reg[96][3]  ( .D(n3120), .CP(clk), .Q(\mem[96][3] ) );
  DFQD1 \mem_reg[96][2]  ( .D(n3119), .CP(clk), .Q(\mem[96][2] ) );
  DFQD1 \mem_reg[96][1]  ( .D(n3118), .CP(clk), .Q(\mem[96][1] ) );
  DFQD1 \mem_reg[96][0]  ( .D(n3117), .CP(clk), .Q(\mem[96][0] ) );
  DFQD1 \mem_reg[97][15]  ( .D(n3116), .CP(clk), .Q(\mem[97][15] ) );
  DFQD1 \mem_reg[97][14]  ( .D(n3115), .CP(clk), .Q(\mem[97][14] ) );
  DFQD1 \mem_reg[97][13]  ( .D(n3114), .CP(clk), .Q(\mem[97][13] ) );
  DFQD1 \mem_reg[97][12]  ( .D(n3113), .CP(clk), .Q(\mem[97][12] ) );
  DFQD1 \mem_reg[97][11]  ( .D(n3112), .CP(clk), .Q(\mem[97][11] ) );
  DFQD1 \mem_reg[97][10]  ( .D(n3111), .CP(clk), .Q(\mem[97][10] ) );
  DFQD1 \mem_reg[97][9]  ( .D(n3110), .CP(clk), .Q(\mem[97][9] ) );
  DFQD1 \mem_reg[97][8]  ( .D(n3109), .CP(clk), .Q(\mem[97][8] ) );
  DFQD1 \mem_reg[97][7]  ( .D(n3108), .CP(clk), .Q(\mem[97][7] ) );
  DFQD1 \mem_reg[97][6]  ( .D(n3107), .CP(clk), .Q(\mem[97][6] ) );
  DFQD1 \mem_reg[97][5]  ( .D(n3106), .CP(clk), .Q(\mem[97][5] ) );
  DFQD1 \mem_reg[97][4]  ( .D(n3105), .CP(clk), .Q(\mem[97][4] ) );
  DFQD1 \mem_reg[97][3]  ( .D(n3104), .CP(clk), .Q(\mem[97][3] ) );
  DFQD1 \mem_reg[97][2]  ( .D(n3103), .CP(clk), .Q(\mem[97][2] ) );
  DFQD1 \mem_reg[97][1]  ( .D(n3102), .CP(clk), .Q(\mem[97][1] ) );
  DFQD1 \mem_reg[97][0]  ( .D(n3101), .CP(clk), .Q(\mem[97][0] ) );
  DFQD1 \mem_reg[98][15]  ( .D(n3100), .CP(clk), .Q(\mem[98][15] ) );
  DFQD1 \mem_reg[98][14]  ( .D(n3099), .CP(clk), .Q(\mem[98][14] ) );
  DFQD1 \mem_reg[98][13]  ( .D(n3098), .CP(clk), .Q(\mem[98][13] ) );
  DFQD1 \mem_reg[98][12]  ( .D(n3097), .CP(clk), .Q(\mem[98][12] ) );
  DFQD1 \mem_reg[98][11]  ( .D(n3096), .CP(clk), .Q(\mem[98][11] ) );
  DFQD1 \mem_reg[98][10]  ( .D(n3095), .CP(clk), .Q(\mem[98][10] ) );
  DFQD1 \mem_reg[98][9]  ( .D(n3094), .CP(clk), .Q(\mem[98][9] ) );
  DFQD1 \mem_reg[98][8]  ( .D(n3093), .CP(clk), .Q(\mem[98][8] ) );
  DFQD1 \mem_reg[98][7]  ( .D(n3092), .CP(clk), .Q(\mem[98][7] ) );
  DFQD1 \mem_reg[98][6]  ( .D(n3091), .CP(clk), .Q(\mem[98][6] ) );
  DFQD1 \mem_reg[98][5]  ( .D(n3090), .CP(clk), .Q(\mem[98][5] ) );
  DFQD1 \mem_reg[98][4]  ( .D(n3089), .CP(clk), .Q(\mem[98][4] ) );
  DFQD1 \mem_reg[98][3]  ( .D(n3088), .CP(clk), .Q(\mem[98][3] ) );
  DFQD1 \mem_reg[98][2]  ( .D(n3087), .CP(clk), .Q(\mem[98][2] ) );
  DFQD1 \mem_reg[98][1]  ( .D(n3086), .CP(clk), .Q(\mem[98][1] ) );
  DFQD1 \mem_reg[98][0]  ( .D(n3085), .CP(clk), .Q(\mem[98][0] ) );
  DFQD1 \mem_reg[99][15]  ( .D(n3084), .CP(clk), .Q(\mem[99][15] ) );
  DFQD1 \mem_reg[99][14]  ( .D(n3083), .CP(clk), .Q(\mem[99][14] ) );
  DFQD1 \mem_reg[99][13]  ( .D(n3082), .CP(clk), .Q(\mem[99][13] ) );
  DFQD1 \mem_reg[99][12]  ( .D(n3081), .CP(clk), .Q(\mem[99][12] ) );
  DFQD1 \mem_reg[99][11]  ( .D(n3080), .CP(clk), .Q(\mem[99][11] ) );
  DFQD1 \mem_reg[99][10]  ( .D(n3079), .CP(clk), .Q(\mem[99][10] ) );
  DFQD1 \mem_reg[99][9]  ( .D(n3078), .CP(clk), .Q(\mem[99][9] ) );
  DFQD1 \mem_reg[99][8]  ( .D(n3077), .CP(clk), .Q(\mem[99][8] ) );
  DFQD1 \mem_reg[99][7]  ( .D(n3076), .CP(clk), .Q(\mem[99][7] ) );
  DFQD1 \mem_reg[99][6]  ( .D(n3075), .CP(clk), .Q(\mem[99][6] ) );
  DFQD1 \mem_reg[99][5]  ( .D(n3074), .CP(clk), .Q(\mem[99][5] ) );
  DFQD1 \mem_reg[99][4]  ( .D(n3073), .CP(clk), .Q(\mem[99][4] ) );
  DFQD1 \mem_reg[99][3]  ( .D(n3072), .CP(clk), .Q(\mem[99][3] ) );
  DFQD1 \mem_reg[99][2]  ( .D(n3071), .CP(clk), .Q(\mem[99][2] ) );
  DFQD1 \mem_reg[99][1]  ( .D(n3070), .CP(clk), .Q(\mem[99][1] ) );
  DFQD1 \mem_reg[99][0]  ( .D(n3069), .CP(clk), .Q(\mem[99][0] ) );
  DFQD1 \mem_reg[100][15]  ( .D(n3068), .CP(clk), .Q(\mem[100][15] ) );
  DFQD1 \mem_reg[100][14]  ( .D(n3067), .CP(clk), .Q(\mem[100][14] ) );
  DFQD1 \mem_reg[100][13]  ( .D(n3066), .CP(clk), .Q(\mem[100][13] ) );
  DFQD1 \mem_reg[100][12]  ( .D(n3065), .CP(clk), .Q(\mem[100][12] ) );
  DFQD1 \mem_reg[100][11]  ( .D(n3064), .CP(clk), .Q(\mem[100][11] ) );
  DFQD1 \mem_reg[100][10]  ( .D(n3063), .CP(clk), .Q(\mem[100][10] ) );
  DFQD1 \mem_reg[100][9]  ( .D(n3062), .CP(clk), .Q(\mem[100][9] ) );
  DFQD1 \mem_reg[100][8]  ( .D(n3061), .CP(clk), .Q(\mem[100][8] ) );
  DFQD1 \mem_reg[100][7]  ( .D(n3060), .CP(clk), .Q(\mem[100][7] ) );
  DFQD1 \mem_reg[100][6]  ( .D(n3059), .CP(clk), .Q(\mem[100][6] ) );
  DFQD1 \mem_reg[100][5]  ( .D(n3058), .CP(clk), .Q(\mem[100][5] ) );
  DFQD1 \mem_reg[100][4]  ( .D(n3057), .CP(clk), .Q(\mem[100][4] ) );
  DFQD1 \mem_reg[100][3]  ( .D(n3056), .CP(clk), .Q(\mem[100][3] ) );
  DFQD1 \mem_reg[100][2]  ( .D(n3055), .CP(clk), .Q(\mem[100][2] ) );
  DFQD1 \mem_reg[100][1]  ( .D(n3054), .CP(clk), .Q(\mem[100][1] ) );
  DFQD1 \mem_reg[100][0]  ( .D(n3053), .CP(clk), .Q(\mem[100][0] ) );
  DFQD1 \mem_reg[101][15]  ( .D(n3052), .CP(clk), .Q(\mem[101][15] ) );
  DFQD1 \mem_reg[101][14]  ( .D(n3051), .CP(clk), .Q(\mem[101][14] ) );
  DFQD1 \mem_reg[101][13]  ( .D(n3050), .CP(clk), .Q(\mem[101][13] ) );
  DFQD1 \mem_reg[101][12]  ( .D(n3049), .CP(clk), .Q(\mem[101][12] ) );
  DFQD1 \mem_reg[101][11]  ( .D(n3048), .CP(clk), .Q(\mem[101][11] ) );
  DFQD1 \mem_reg[101][10]  ( .D(n3047), .CP(clk), .Q(\mem[101][10] ) );
  DFQD1 \mem_reg[101][9]  ( .D(n3046), .CP(clk), .Q(\mem[101][9] ) );
  DFQD1 \mem_reg[101][8]  ( .D(n3045), .CP(clk), .Q(\mem[101][8] ) );
  DFQD1 \mem_reg[101][7]  ( .D(n3044), .CP(clk), .Q(\mem[101][7] ) );
  DFQD1 \mem_reg[101][6]  ( .D(n3043), .CP(clk), .Q(\mem[101][6] ) );
  DFQD1 \mem_reg[101][5]  ( .D(n3042), .CP(clk), .Q(\mem[101][5] ) );
  DFQD1 \mem_reg[101][4]  ( .D(n3041), .CP(clk), .Q(\mem[101][4] ) );
  DFQD1 \mem_reg[101][3]  ( .D(n3040), .CP(clk), .Q(\mem[101][3] ) );
  DFQD1 \mem_reg[101][2]  ( .D(n3039), .CP(clk), .Q(\mem[101][2] ) );
  DFQD1 \mem_reg[101][1]  ( .D(n3038), .CP(clk), .Q(\mem[101][1] ) );
  DFQD1 \mem_reg[101][0]  ( .D(n3037), .CP(clk), .Q(\mem[101][0] ) );
  DFQD1 \mem_reg[102][15]  ( .D(n3036), .CP(clk), .Q(\mem[102][15] ) );
  DFQD1 \mem_reg[102][14]  ( .D(n3035), .CP(clk), .Q(\mem[102][14] ) );
  DFQD1 \mem_reg[102][13]  ( .D(n3034), .CP(clk), .Q(\mem[102][13] ) );
  DFQD1 \mem_reg[102][12]  ( .D(n3033), .CP(clk), .Q(\mem[102][12] ) );
  DFQD1 \mem_reg[102][11]  ( .D(n3032), .CP(clk), .Q(\mem[102][11] ) );
  DFQD1 \mem_reg[102][10]  ( .D(n3031), .CP(clk), .Q(\mem[102][10] ) );
  DFQD1 \mem_reg[102][9]  ( .D(n3030), .CP(clk), .Q(\mem[102][9] ) );
  DFQD1 \mem_reg[102][8]  ( .D(n3029), .CP(clk), .Q(\mem[102][8] ) );
  DFQD1 \mem_reg[102][7]  ( .D(n3028), .CP(clk), .Q(\mem[102][7] ) );
  DFQD1 \mem_reg[102][6]  ( .D(n3027), .CP(clk), .Q(\mem[102][6] ) );
  DFQD1 \mem_reg[102][5]  ( .D(n3026), .CP(clk), .Q(\mem[102][5] ) );
  DFQD1 \mem_reg[102][4]  ( .D(n3025), .CP(clk), .Q(\mem[102][4] ) );
  DFQD1 \mem_reg[102][3]  ( .D(n3024), .CP(clk), .Q(\mem[102][3] ) );
  DFQD1 \mem_reg[102][2]  ( .D(n3023), .CP(clk), .Q(\mem[102][2] ) );
  DFQD1 \mem_reg[102][1]  ( .D(n3022), .CP(clk), .Q(\mem[102][1] ) );
  DFQD1 \mem_reg[102][0]  ( .D(n3021), .CP(clk), .Q(\mem[102][0] ) );
  DFQD1 \mem_reg[103][15]  ( .D(n3020), .CP(clk), .Q(\mem[103][15] ) );
  DFQD1 \mem_reg[103][14]  ( .D(n3019), .CP(clk), .Q(\mem[103][14] ) );
  DFQD1 \mem_reg[103][13]  ( .D(n3018), .CP(clk), .Q(\mem[103][13] ) );
  DFQD1 \mem_reg[103][12]  ( .D(n3017), .CP(clk), .Q(\mem[103][12] ) );
  DFQD1 \mem_reg[103][11]  ( .D(n3016), .CP(clk), .Q(\mem[103][11] ) );
  DFQD1 \mem_reg[103][10]  ( .D(n3015), .CP(clk), .Q(\mem[103][10] ) );
  DFQD1 \mem_reg[103][9]  ( .D(n3014), .CP(clk), .Q(\mem[103][9] ) );
  DFQD1 \mem_reg[103][8]  ( .D(n3013), .CP(clk), .Q(\mem[103][8] ) );
  DFQD1 \mem_reg[103][7]  ( .D(n3012), .CP(clk), .Q(\mem[103][7] ) );
  DFQD1 \mem_reg[103][6]  ( .D(n3011), .CP(clk), .Q(\mem[103][6] ) );
  DFQD1 \mem_reg[103][5]  ( .D(n3010), .CP(clk), .Q(\mem[103][5] ) );
  DFQD1 \mem_reg[103][4]  ( .D(n3009), .CP(clk), .Q(\mem[103][4] ) );
  DFQD1 \mem_reg[103][3]  ( .D(n3008), .CP(clk), .Q(\mem[103][3] ) );
  DFQD1 \mem_reg[103][2]  ( .D(n3007), .CP(clk), .Q(\mem[103][2] ) );
  DFQD1 \mem_reg[103][1]  ( .D(n3006), .CP(clk), .Q(\mem[103][1] ) );
  DFQD1 \mem_reg[103][0]  ( .D(n3005), .CP(clk), .Q(\mem[103][0] ) );
  DFQD1 \mem_reg[104][15]  ( .D(n3004), .CP(clk), .Q(\mem[104][15] ) );
  DFQD1 \mem_reg[104][14]  ( .D(n3003), .CP(clk), .Q(\mem[104][14] ) );
  DFQD1 \mem_reg[104][13]  ( .D(n3002), .CP(clk), .Q(\mem[104][13] ) );
  DFQD1 \mem_reg[104][12]  ( .D(n3001), .CP(clk), .Q(\mem[104][12] ) );
  DFQD1 \mem_reg[104][11]  ( .D(n3000), .CP(clk), .Q(\mem[104][11] ) );
  DFQD1 \mem_reg[104][10]  ( .D(n2999), .CP(clk), .Q(\mem[104][10] ) );
  DFQD1 \mem_reg[104][9]  ( .D(n2998), .CP(clk), .Q(\mem[104][9] ) );
  DFQD1 \mem_reg[104][8]  ( .D(n2997), .CP(clk), .Q(\mem[104][8] ) );
  DFQD1 \mem_reg[104][7]  ( .D(n2996), .CP(clk), .Q(\mem[104][7] ) );
  DFQD1 \mem_reg[104][6]  ( .D(n2995), .CP(clk), .Q(\mem[104][6] ) );
  DFQD1 \mem_reg[104][5]  ( .D(n2994), .CP(clk), .Q(\mem[104][5] ) );
  DFQD1 \mem_reg[104][4]  ( .D(n2993), .CP(clk), .Q(\mem[104][4] ) );
  DFQD1 \mem_reg[104][3]  ( .D(n2992), .CP(clk), .Q(\mem[104][3] ) );
  DFQD1 \mem_reg[104][2]  ( .D(n2991), .CP(clk), .Q(\mem[104][2] ) );
  DFQD1 \mem_reg[104][1]  ( .D(n2990), .CP(clk), .Q(\mem[104][1] ) );
  DFQD1 \mem_reg[104][0]  ( .D(n2989), .CP(clk), .Q(\mem[104][0] ) );
  DFQD1 \mem_reg[105][15]  ( .D(n2988), .CP(clk), .Q(\mem[105][15] ) );
  DFQD1 \mem_reg[105][14]  ( .D(n2987), .CP(clk), .Q(\mem[105][14] ) );
  DFQD1 \mem_reg[105][13]  ( .D(n2986), .CP(clk), .Q(\mem[105][13] ) );
  DFQD1 \mem_reg[105][12]  ( .D(n2985), .CP(clk), .Q(\mem[105][12] ) );
  DFQD1 \mem_reg[105][11]  ( .D(n2984), .CP(clk), .Q(\mem[105][11] ) );
  DFQD1 \mem_reg[105][10]  ( .D(n2983), .CP(clk), .Q(\mem[105][10] ) );
  DFQD1 \mem_reg[105][9]  ( .D(n2982), .CP(clk), .Q(\mem[105][9] ) );
  DFQD1 \mem_reg[105][8]  ( .D(n2981), .CP(clk), .Q(\mem[105][8] ) );
  DFQD1 \mem_reg[105][7]  ( .D(n2980), .CP(clk), .Q(\mem[105][7] ) );
  DFQD1 \mem_reg[105][6]  ( .D(n2979), .CP(clk), .Q(\mem[105][6] ) );
  DFQD1 \mem_reg[105][5]  ( .D(n2978), .CP(clk), .Q(\mem[105][5] ) );
  DFQD1 \mem_reg[105][4]  ( .D(n2977), .CP(clk), .Q(\mem[105][4] ) );
  DFQD1 \mem_reg[105][3]  ( .D(n2976), .CP(clk), .Q(\mem[105][3] ) );
  DFQD1 \mem_reg[105][2]  ( .D(n2975), .CP(clk), .Q(\mem[105][2] ) );
  DFQD1 \mem_reg[105][1]  ( .D(n2974), .CP(clk), .Q(\mem[105][1] ) );
  DFQD1 \mem_reg[105][0]  ( .D(n2973), .CP(clk), .Q(\mem[105][0] ) );
  DFQD1 \mem_reg[106][15]  ( .D(n2972), .CP(clk), .Q(\mem[106][15] ) );
  DFQD1 \mem_reg[106][14]  ( .D(n2971), .CP(clk), .Q(\mem[106][14] ) );
  DFQD1 \mem_reg[106][13]  ( .D(n2970), .CP(clk), .Q(\mem[106][13] ) );
  DFQD1 \mem_reg[106][12]  ( .D(n2969), .CP(clk), .Q(\mem[106][12] ) );
  DFQD1 \mem_reg[106][11]  ( .D(n2968), .CP(clk), .Q(\mem[106][11] ) );
  DFQD1 \mem_reg[106][10]  ( .D(n2967), .CP(clk), .Q(\mem[106][10] ) );
  DFQD1 \mem_reg[106][9]  ( .D(n2966), .CP(clk), .Q(\mem[106][9] ) );
  DFQD1 \mem_reg[106][8]  ( .D(n2965), .CP(clk), .Q(\mem[106][8] ) );
  DFQD1 \mem_reg[106][7]  ( .D(n2964), .CP(clk), .Q(\mem[106][7] ) );
  DFQD1 \mem_reg[106][6]  ( .D(n2963), .CP(clk), .Q(\mem[106][6] ) );
  DFQD1 \mem_reg[106][5]  ( .D(n2962), .CP(clk), .Q(\mem[106][5] ) );
  DFQD1 \mem_reg[106][4]  ( .D(n2961), .CP(clk), .Q(\mem[106][4] ) );
  DFQD1 \mem_reg[106][3]  ( .D(n2960), .CP(clk), .Q(\mem[106][3] ) );
  DFQD1 \mem_reg[106][2]  ( .D(n2959), .CP(clk), .Q(\mem[106][2] ) );
  DFQD1 \mem_reg[106][1]  ( .D(n2958), .CP(clk), .Q(\mem[106][1] ) );
  DFQD1 \mem_reg[106][0]  ( .D(n2957), .CP(clk), .Q(\mem[106][0] ) );
  DFQD1 \mem_reg[107][15]  ( .D(n2956), .CP(clk), .Q(\mem[107][15] ) );
  DFQD1 \mem_reg[107][14]  ( .D(n2955), .CP(clk), .Q(\mem[107][14] ) );
  DFQD1 \mem_reg[107][13]  ( .D(n2954), .CP(clk), .Q(\mem[107][13] ) );
  DFQD1 \mem_reg[107][12]  ( .D(n2953), .CP(clk), .Q(\mem[107][12] ) );
  DFQD1 \mem_reg[107][11]  ( .D(n2952), .CP(clk), .Q(\mem[107][11] ) );
  DFQD1 \mem_reg[107][10]  ( .D(n2951), .CP(clk), .Q(\mem[107][10] ) );
  DFQD1 \mem_reg[107][9]  ( .D(n2950), .CP(clk), .Q(\mem[107][9] ) );
  DFQD1 \mem_reg[107][8]  ( .D(n2949), .CP(clk), .Q(\mem[107][8] ) );
  DFQD1 \mem_reg[107][7]  ( .D(n2948), .CP(clk), .Q(\mem[107][7] ) );
  DFQD1 \mem_reg[107][6]  ( .D(n2947), .CP(clk), .Q(\mem[107][6] ) );
  DFQD1 \mem_reg[107][5]  ( .D(n2946), .CP(clk), .Q(\mem[107][5] ) );
  DFQD1 \mem_reg[107][4]  ( .D(n2945), .CP(clk), .Q(\mem[107][4] ) );
  DFQD1 \mem_reg[107][3]  ( .D(n2944), .CP(clk), .Q(\mem[107][3] ) );
  DFQD1 \mem_reg[107][2]  ( .D(n2943), .CP(clk), .Q(\mem[107][2] ) );
  DFQD1 \mem_reg[107][1]  ( .D(n2942), .CP(clk), .Q(\mem[107][1] ) );
  DFQD1 \mem_reg[107][0]  ( .D(n2941), .CP(clk), .Q(\mem[107][0] ) );
  DFQD1 \mem_reg[108][15]  ( .D(n2940), .CP(clk), .Q(\mem[108][15] ) );
  DFQD1 \mem_reg[108][14]  ( .D(n2939), .CP(clk), .Q(\mem[108][14] ) );
  DFQD1 \mem_reg[108][13]  ( .D(n2938), .CP(clk), .Q(\mem[108][13] ) );
  DFQD1 \mem_reg[108][12]  ( .D(n2937), .CP(clk), .Q(\mem[108][12] ) );
  DFQD1 \mem_reg[108][11]  ( .D(n2936), .CP(clk), .Q(\mem[108][11] ) );
  DFQD1 \mem_reg[108][10]  ( .D(n2935), .CP(clk), .Q(\mem[108][10] ) );
  DFQD1 \mem_reg[108][9]  ( .D(n2934), .CP(clk), .Q(\mem[108][9] ) );
  DFQD1 \mem_reg[108][8]  ( .D(n2933), .CP(clk), .Q(\mem[108][8] ) );
  DFQD1 \mem_reg[108][7]  ( .D(n2932), .CP(clk), .Q(\mem[108][7] ) );
  DFQD1 \mem_reg[108][6]  ( .D(n2931), .CP(clk), .Q(\mem[108][6] ) );
  DFQD1 \mem_reg[108][5]  ( .D(n2930), .CP(clk), .Q(\mem[108][5] ) );
  DFQD1 \mem_reg[108][4]  ( .D(n2929), .CP(clk), .Q(\mem[108][4] ) );
  DFQD1 \mem_reg[108][3]  ( .D(n2928), .CP(clk), .Q(\mem[108][3] ) );
  DFQD1 \mem_reg[108][2]  ( .D(n2927), .CP(clk), .Q(\mem[108][2] ) );
  DFQD1 \mem_reg[108][1]  ( .D(n2926), .CP(clk), .Q(\mem[108][1] ) );
  DFQD1 \mem_reg[108][0]  ( .D(n2925), .CP(clk), .Q(\mem[108][0] ) );
  DFQD1 \mem_reg[109][15]  ( .D(n2924), .CP(clk), .Q(\mem[109][15] ) );
  DFQD1 \mem_reg[109][14]  ( .D(n2923), .CP(clk), .Q(\mem[109][14] ) );
  DFQD1 \mem_reg[109][13]  ( .D(n2922), .CP(clk), .Q(\mem[109][13] ) );
  DFQD1 \mem_reg[109][12]  ( .D(n2921), .CP(clk), .Q(\mem[109][12] ) );
  DFQD1 \mem_reg[109][11]  ( .D(n2920), .CP(clk), .Q(\mem[109][11] ) );
  DFQD1 \mem_reg[109][10]  ( .D(n2919), .CP(clk), .Q(\mem[109][10] ) );
  DFQD1 \mem_reg[109][9]  ( .D(n2918), .CP(clk), .Q(\mem[109][9] ) );
  DFQD1 \mem_reg[109][8]  ( .D(n2917), .CP(clk), .Q(\mem[109][8] ) );
  DFQD1 \mem_reg[109][7]  ( .D(n2916), .CP(clk), .Q(\mem[109][7] ) );
  DFQD1 \mem_reg[109][6]  ( .D(n2915), .CP(clk), .Q(\mem[109][6] ) );
  DFQD1 \mem_reg[109][5]  ( .D(n2914), .CP(clk), .Q(\mem[109][5] ) );
  DFQD1 \mem_reg[109][4]  ( .D(n2913), .CP(clk), .Q(\mem[109][4] ) );
  DFQD1 \mem_reg[109][3]  ( .D(n2912), .CP(clk), .Q(\mem[109][3] ) );
  DFQD1 \mem_reg[109][2]  ( .D(n2911), .CP(clk), .Q(\mem[109][2] ) );
  DFQD1 \mem_reg[109][1]  ( .D(n2910), .CP(clk), .Q(\mem[109][1] ) );
  DFQD1 \mem_reg[109][0]  ( .D(n2909), .CP(clk), .Q(\mem[109][0] ) );
  DFQD1 \mem_reg[110][15]  ( .D(n2908), .CP(clk), .Q(\mem[110][15] ) );
  DFQD1 \mem_reg[110][14]  ( .D(n2907), .CP(clk), .Q(\mem[110][14] ) );
  DFQD1 \mem_reg[110][13]  ( .D(n2906), .CP(clk), .Q(\mem[110][13] ) );
  DFQD1 \mem_reg[110][12]  ( .D(n2905), .CP(clk), .Q(\mem[110][12] ) );
  DFQD1 \mem_reg[110][11]  ( .D(n2904), .CP(clk), .Q(\mem[110][11] ) );
  DFQD1 \mem_reg[110][10]  ( .D(n2903), .CP(clk), .Q(\mem[110][10] ) );
  DFQD1 \mem_reg[110][9]  ( .D(n2902), .CP(clk), .Q(\mem[110][9] ) );
  DFQD1 \mem_reg[110][8]  ( .D(n2901), .CP(clk), .Q(\mem[110][8] ) );
  DFQD1 \mem_reg[110][7]  ( .D(n2900), .CP(clk), .Q(\mem[110][7] ) );
  DFQD1 \mem_reg[110][6]  ( .D(n2899), .CP(clk), .Q(\mem[110][6] ) );
  DFQD1 \mem_reg[110][5]  ( .D(n2898), .CP(clk), .Q(\mem[110][5] ) );
  DFQD1 \mem_reg[110][4]  ( .D(n2897), .CP(clk), .Q(\mem[110][4] ) );
  DFQD1 \mem_reg[110][3]  ( .D(n2896), .CP(clk), .Q(\mem[110][3] ) );
  DFQD1 \mem_reg[110][2]  ( .D(n2895), .CP(clk), .Q(\mem[110][2] ) );
  DFQD1 \mem_reg[110][1]  ( .D(n2894), .CP(clk), .Q(\mem[110][1] ) );
  DFQD1 \mem_reg[110][0]  ( .D(n2893), .CP(clk), .Q(\mem[110][0] ) );
  DFQD1 \mem_reg[111][15]  ( .D(n2892), .CP(clk), .Q(\mem[111][15] ) );
  DFQD1 \mem_reg[111][14]  ( .D(n2891), .CP(clk), .Q(\mem[111][14] ) );
  DFQD1 \mem_reg[111][13]  ( .D(n2890), .CP(clk), .Q(\mem[111][13] ) );
  DFQD1 \mem_reg[111][12]  ( .D(n2889), .CP(clk), .Q(\mem[111][12] ) );
  DFQD1 \mem_reg[111][11]  ( .D(n2888), .CP(clk), .Q(\mem[111][11] ) );
  DFQD1 \mem_reg[111][10]  ( .D(n2887), .CP(clk), .Q(\mem[111][10] ) );
  DFQD1 \mem_reg[111][9]  ( .D(n2886), .CP(clk), .Q(\mem[111][9] ) );
  DFQD1 \mem_reg[111][8]  ( .D(n2885), .CP(clk), .Q(\mem[111][8] ) );
  DFQD1 \mem_reg[111][7]  ( .D(n2884), .CP(clk), .Q(\mem[111][7] ) );
  DFQD1 \mem_reg[111][6]  ( .D(n2883), .CP(clk), .Q(\mem[111][6] ) );
  DFQD1 \mem_reg[111][5]  ( .D(n2882), .CP(clk), .Q(\mem[111][5] ) );
  DFQD1 \mem_reg[111][4]  ( .D(n2881), .CP(clk), .Q(\mem[111][4] ) );
  DFQD1 \mem_reg[111][3]  ( .D(n2880), .CP(clk), .Q(\mem[111][3] ) );
  DFQD1 \mem_reg[111][2]  ( .D(n2879), .CP(clk), .Q(\mem[111][2] ) );
  DFQD1 \mem_reg[111][1]  ( .D(n2878), .CP(clk), .Q(\mem[111][1] ) );
  DFQD1 \mem_reg[111][0]  ( .D(n2877), .CP(clk), .Q(\mem[111][0] ) );
  DFQD1 \mem_reg[112][15]  ( .D(n2876), .CP(clk), .Q(\mem[112][15] ) );
  DFQD1 \mem_reg[112][14]  ( .D(n2875), .CP(clk), .Q(\mem[112][14] ) );
  DFQD1 \mem_reg[112][13]  ( .D(n2874), .CP(clk), .Q(\mem[112][13] ) );
  DFQD1 \mem_reg[112][12]  ( .D(n2873), .CP(clk), .Q(\mem[112][12] ) );
  DFQD1 \mem_reg[112][11]  ( .D(n2872), .CP(clk), .Q(\mem[112][11] ) );
  DFQD1 \mem_reg[112][10]  ( .D(n2871), .CP(clk), .Q(\mem[112][10] ) );
  DFQD1 \mem_reg[112][9]  ( .D(n2870), .CP(clk), .Q(\mem[112][9] ) );
  DFQD1 \mem_reg[112][8]  ( .D(n2869), .CP(clk), .Q(\mem[112][8] ) );
  DFQD1 \mem_reg[112][7]  ( .D(n2868), .CP(clk), .Q(\mem[112][7] ) );
  DFQD1 \mem_reg[112][6]  ( .D(n2867), .CP(clk), .Q(\mem[112][6] ) );
  DFQD1 \mem_reg[112][5]  ( .D(n2866), .CP(clk), .Q(\mem[112][5] ) );
  DFQD1 \mem_reg[112][4]  ( .D(n2865), .CP(clk), .Q(\mem[112][4] ) );
  DFQD1 \mem_reg[112][3]  ( .D(n2864), .CP(clk), .Q(\mem[112][3] ) );
  DFQD1 \mem_reg[112][2]  ( .D(n2863), .CP(clk), .Q(\mem[112][2] ) );
  DFQD1 \mem_reg[112][1]  ( .D(n2862), .CP(clk), .Q(\mem[112][1] ) );
  DFQD1 \mem_reg[112][0]  ( .D(n2861), .CP(clk), .Q(\mem[112][0] ) );
  DFQD1 \mem_reg[113][15]  ( .D(n2860), .CP(clk), .Q(\mem[113][15] ) );
  DFQD1 \mem_reg[113][14]  ( .D(n2859), .CP(clk), .Q(\mem[113][14] ) );
  DFQD1 \mem_reg[113][13]  ( .D(n2858), .CP(clk), .Q(\mem[113][13] ) );
  DFQD1 \mem_reg[113][12]  ( .D(n2857), .CP(clk), .Q(\mem[113][12] ) );
  DFQD1 \mem_reg[113][11]  ( .D(n2856), .CP(clk), .Q(\mem[113][11] ) );
  DFQD1 \mem_reg[113][10]  ( .D(n2855), .CP(clk), .Q(\mem[113][10] ) );
  DFQD1 \mem_reg[113][9]  ( .D(n2854), .CP(clk), .Q(\mem[113][9] ) );
  DFQD1 \mem_reg[113][8]  ( .D(n2853), .CP(clk), .Q(\mem[113][8] ) );
  DFQD1 \mem_reg[113][7]  ( .D(n2852), .CP(clk), .Q(\mem[113][7] ) );
  DFQD1 \mem_reg[113][6]  ( .D(n2851), .CP(clk), .Q(\mem[113][6] ) );
  DFQD1 \mem_reg[113][5]  ( .D(n2850), .CP(clk), .Q(\mem[113][5] ) );
  DFQD1 \mem_reg[113][4]  ( .D(n2849), .CP(clk), .Q(\mem[113][4] ) );
  DFQD1 \mem_reg[113][3]  ( .D(n2848), .CP(clk), .Q(\mem[113][3] ) );
  DFQD1 \mem_reg[113][2]  ( .D(n2847), .CP(clk), .Q(\mem[113][2] ) );
  DFQD1 \mem_reg[113][1]  ( .D(n2846), .CP(clk), .Q(\mem[113][1] ) );
  DFQD1 \mem_reg[113][0]  ( .D(n2845), .CP(clk), .Q(\mem[113][0] ) );
  DFQD1 \mem_reg[114][15]  ( .D(n2844), .CP(clk), .Q(\mem[114][15] ) );
  DFQD1 \mem_reg[114][14]  ( .D(n2843), .CP(clk), .Q(\mem[114][14] ) );
  DFQD1 \mem_reg[114][13]  ( .D(n2842), .CP(clk), .Q(\mem[114][13] ) );
  DFQD1 \mem_reg[114][12]  ( .D(n2841), .CP(clk), .Q(\mem[114][12] ) );
  DFQD1 \mem_reg[114][11]  ( .D(n2840), .CP(clk), .Q(\mem[114][11] ) );
  DFQD1 \mem_reg[114][10]  ( .D(n2839), .CP(clk), .Q(\mem[114][10] ) );
  DFQD1 \mem_reg[114][9]  ( .D(n2838), .CP(clk), .Q(\mem[114][9] ) );
  DFQD1 \mem_reg[114][8]  ( .D(n2837), .CP(clk), .Q(\mem[114][8] ) );
  DFQD1 \mem_reg[114][7]  ( .D(n2836), .CP(clk), .Q(\mem[114][7] ) );
  DFQD1 \mem_reg[114][6]  ( .D(n2835), .CP(clk), .Q(\mem[114][6] ) );
  DFQD1 \mem_reg[114][5]  ( .D(n2834), .CP(clk), .Q(\mem[114][5] ) );
  DFQD1 \mem_reg[114][4]  ( .D(n2833), .CP(clk), .Q(\mem[114][4] ) );
  DFQD1 \mem_reg[114][3]  ( .D(n2832), .CP(clk), .Q(\mem[114][3] ) );
  DFQD1 \mem_reg[114][2]  ( .D(n2831), .CP(clk), .Q(\mem[114][2] ) );
  DFQD1 \mem_reg[114][1]  ( .D(n2830), .CP(clk), .Q(\mem[114][1] ) );
  DFQD1 \mem_reg[114][0]  ( .D(n2829), .CP(clk), .Q(\mem[114][0] ) );
  DFQD1 \mem_reg[115][15]  ( .D(n2828), .CP(clk), .Q(\mem[115][15] ) );
  DFQD1 \mem_reg[115][14]  ( .D(n2827), .CP(clk), .Q(\mem[115][14] ) );
  DFQD1 \mem_reg[115][13]  ( .D(n2826), .CP(clk), .Q(\mem[115][13] ) );
  DFQD1 \mem_reg[115][12]  ( .D(n2825), .CP(clk), .Q(\mem[115][12] ) );
  DFQD1 \mem_reg[115][11]  ( .D(n2824), .CP(clk), .Q(\mem[115][11] ) );
  DFQD1 \mem_reg[115][10]  ( .D(n2823), .CP(clk), .Q(\mem[115][10] ) );
  DFQD1 \mem_reg[115][9]  ( .D(n2822), .CP(clk), .Q(\mem[115][9] ) );
  DFQD1 \mem_reg[115][8]  ( .D(n2821), .CP(clk), .Q(\mem[115][8] ) );
  DFQD1 \mem_reg[115][7]  ( .D(n2820), .CP(clk), .Q(\mem[115][7] ) );
  DFQD1 \mem_reg[115][6]  ( .D(n2819), .CP(clk), .Q(\mem[115][6] ) );
  DFQD1 \mem_reg[115][5]  ( .D(n2818), .CP(clk), .Q(\mem[115][5] ) );
  DFQD1 \mem_reg[115][4]  ( .D(n2817), .CP(clk), .Q(\mem[115][4] ) );
  DFQD1 \mem_reg[115][3]  ( .D(n2816), .CP(clk), .Q(\mem[115][3] ) );
  DFQD1 \mem_reg[115][2]  ( .D(n2815), .CP(clk), .Q(\mem[115][2] ) );
  DFQD1 \mem_reg[115][1]  ( .D(n2814), .CP(clk), .Q(\mem[115][1] ) );
  DFQD1 \mem_reg[115][0]  ( .D(n2813), .CP(clk), .Q(\mem[115][0] ) );
  DFQD1 \mem_reg[116][15]  ( .D(n2812), .CP(clk), .Q(\mem[116][15] ) );
  DFQD1 \mem_reg[116][14]  ( .D(n2811), .CP(clk), .Q(\mem[116][14] ) );
  DFQD1 \mem_reg[116][13]  ( .D(n2810), .CP(clk), .Q(\mem[116][13] ) );
  DFQD1 \mem_reg[116][12]  ( .D(n2809), .CP(clk), .Q(\mem[116][12] ) );
  DFQD1 \mem_reg[116][11]  ( .D(n2808), .CP(clk), .Q(\mem[116][11] ) );
  DFQD1 \mem_reg[116][10]  ( .D(n2807), .CP(clk), .Q(\mem[116][10] ) );
  DFQD1 \mem_reg[116][9]  ( .D(n2806), .CP(clk), .Q(\mem[116][9] ) );
  DFQD1 \mem_reg[116][8]  ( .D(n2805), .CP(clk), .Q(\mem[116][8] ) );
  DFQD1 \mem_reg[116][7]  ( .D(n2804), .CP(clk), .Q(\mem[116][7] ) );
  DFQD1 \mem_reg[116][6]  ( .D(n2803), .CP(clk), .Q(\mem[116][6] ) );
  DFQD1 \mem_reg[116][5]  ( .D(n2802), .CP(clk), .Q(\mem[116][5] ) );
  DFQD1 \mem_reg[116][4]  ( .D(n2801), .CP(clk), .Q(\mem[116][4] ) );
  DFQD1 \mem_reg[116][3]  ( .D(n2800), .CP(clk), .Q(\mem[116][3] ) );
  DFQD1 \mem_reg[116][2]  ( .D(n2799), .CP(clk), .Q(\mem[116][2] ) );
  DFQD1 \mem_reg[116][1]  ( .D(n2798), .CP(clk), .Q(\mem[116][1] ) );
  DFQD1 \mem_reg[116][0]  ( .D(n2797), .CP(clk), .Q(\mem[116][0] ) );
  DFQD1 \mem_reg[117][15]  ( .D(n2796), .CP(clk), .Q(\mem[117][15] ) );
  DFQD1 \mem_reg[117][14]  ( .D(n2795), .CP(clk), .Q(\mem[117][14] ) );
  DFQD1 \mem_reg[117][13]  ( .D(n2794), .CP(clk), .Q(\mem[117][13] ) );
  DFQD1 \mem_reg[117][12]  ( .D(n2793), .CP(clk), .Q(\mem[117][12] ) );
  DFQD1 \mem_reg[117][11]  ( .D(n2792), .CP(clk), .Q(\mem[117][11] ) );
  DFQD1 \mem_reg[117][10]  ( .D(n2791), .CP(clk), .Q(\mem[117][10] ) );
  DFQD1 \mem_reg[117][9]  ( .D(n2790), .CP(clk), .Q(\mem[117][9] ) );
  DFQD1 \mem_reg[117][8]  ( .D(n2789), .CP(clk), .Q(\mem[117][8] ) );
  DFQD1 \mem_reg[117][7]  ( .D(n2788), .CP(clk), .Q(\mem[117][7] ) );
  DFQD1 \mem_reg[117][6]  ( .D(n2787), .CP(clk), .Q(\mem[117][6] ) );
  DFQD1 \mem_reg[117][5]  ( .D(n2786), .CP(clk), .Q(\mem[117][5] ) );
  DFQD1 \mem_reg[117][4]  ( .D(n2785), .CP(clk), .Q(\mem[117][4] ) );
  DFQD1 \mem_reg[117][3]  ( .D(n2784), .CP(clk), .Q(\mem[117][3] ) );
  DFQD1 \mem_reg[117][2]  ( .D(n2783), .CP(clk), .Q(\mem[117][2] ) );
  DFQD1 \mem_reg[117][1]  ( .D(n2782), .CP(clk), .Q(\mem[117][1] ) );
  DFQD1 \mem_reg[117][0]  ( .D(n2781), .CP(clk), .Q(\mem[117][0] ) );
  DFQD1 \mem_reg[118][15]  ( .D(n2780), .CP(clk), .Q(\mem[118][15] ) );
  DFQD1 \mem_reg[118][14]  ( .D(n2779), .CP(clk), .Q(\mem[118][14] ) );
  DFQD1 \mem_reg[118][13]  ( .D(n2778), .CP(clk), .Q(\mem[118][13] ) );
  DFQD1 \mem_reg[118][12]  ( .D(n2777), .CP(clk), .Q(\mem[118][12] ) );
  DFQD1 \mem_reg[118][11]  ( .D(n2776), .CP(clk), .Q(\mem[118][11] ) );
  DFQD1 \mem_reg[118][10]  ( .D(n2775), .CP(clk), .Q(\mem[118][10] ) );
  DFQD1 \mem_reg[118][9]  ( .D(n2774), .CP(clk), .Q(\mem[118][9] ) );
  DFQD1 \mem_reg[118][8]  ( .D(n2773), .CP(clk), .Q(\mem[118][8] ) );
  DFQD1 \mem_reg[118][7]  ( .D(n2772), .CP(clk), .Q(\mem[118][7] ) );
  DFQD1 \mem_reg[118][6]  ( .D(n2771), .CP(clk), .Q(\mem[118][6] ) );
  DFQD1 \mem_reg[118][5]  ( .D(n2770), .CP(clk), .Q(\mem[118][5] ) );
  DFQD1 \mem_reg[118][4]  ( .D(n2769), .CP(clk), .Q(\mem[118][4] ) );
  DFQD1 \mem_reg[118][3]  ( .D(n2768), .CP(clk), .Q(\mem[118][3] ) );
  DFQD1 \mem_reg[118][2]  ( .D(n2767), .CP(clk), .Q(\mem[118][2] ) );
  DFQD1 \mem_reg[118][1]  ( .D(n2766), .CP(clk), .Q(\mem[118][1] ) );
  DFQD1 \mem_reg[118][0]  ( .D(n2765), .CP(clk), .Q(\mem[118][0] ) );
  DFQD1 \mem_reg[119][15]  ( .D(n2764), .CP(clk), .Q(\mem[119][15] ) );
  DFQD1 \mem_reg[119][14]  ( .D(n2763), .CP(clk), .Q(\mem[119][14] ) );
  DFQD1 \mem_reg[119][13]  ( .D(n2762), .CP(clk), .Q(\mem[119][13] ) );
  DFQD1 \mem_reg[119][12]  ( .D(n2761), .CP(clk), .Q(\mem[119][12] ) );
  DFQD1 \mem_reg[119][11]  ( .D(n2760), .CP(clk), .Q(\mem[119][11] ) );
  DFQD1 \mem_reg[119][10]  ( .D(n2759), .CP(clk), .Q(\mem[119][10] ) );
  DFQD1 \mem_reg[119][9]  ( .D(n2758), .CP(clk), .Q(\mem[119][9] ) );
  DFQD1 \mem_reg[119][8]  ( .D(n2757), .CP(clk), .Q(\mem[119][8] ) );
  DFQD1 \mem_reg[119][7]  ( .D(n2756), .CP(clk), .Q(\mem[119][7] ) );
  DFQD1 \mem_reg[119][6]  ( .D(n2755), .CP(clk), .Q(\mem[119][6] ) );
  DFQD1 \mem_reg[119][5]  ( .D(n2754), .CP(clk), .Q(\mem[119][5] ) );
  DFQD1 \mem_reg[119][4]  ( .D(n2753), .CP(clk), .Q(\mem[119][4] ) );
  DFQD1 \mem_reg[119][3]  ( .D(n2752), .CP(clk), .Q(\mem[119][3] ) );
  DFQD1 \mem_reg[119][2]  ( .D(n2751), .CP(clk), .Q(\mem[119][2] ) );
  DFQD1 \mem_reg[119][1]  ( .D(n2750), .CP(clk), .Q(\mem[119][1] ) );
  DFQD1 \mem_reg[119][0]  ( .D(n2749), .CP(clk), .Q(\mem[119][0] ) );
  DFQD1 \mem_reg[120][15]  ( .D(n2748), .CP(clk), .Q(\mem[120][15] ) );
  DFQD1 \mem_reg[120][14]  ( .D(n2747), .CP(clk), .Q(\mem[120][14] ) );
  DFQD1 \mem_reg[120][13]  ( .D(n2746), .CP(clk), .Q(\mem[120][13] ) );
  DFQD1 \mem_reg[120][12]  ( .D(n2745), .CP(clk), .Q(\mem[120][12] ) );
  DFQD1 \mem_reg[120][11]  ( .D(n2744), .CP(clk), .Q(\mem[120][11] ) );
  DFQD1 \mem_reg[120][10]  ( .D(n2743), .CP(clk), .Q(\mem[120][10] ) );
  DFQD1 \mem_reg[120][9]  ( .D(n2742), .CP(clk), .Q(\mem[120][9] ) );
  DFQD1 \mem_reg[120][8]  ( .D(n2741), .CP(clk), .Q(\mem[120][8] ) );
  DFQD1 \mem_reg[120][7]  ( .D(n2740), .CP(clk), .Q(\mem[120][7] ) );
  DFQD1 \mem_reg[120][6]  ( .D(n2739), .CP(clk), .Q(\mem[120][6] ) );
  DFQD1 \mem_reg[120][5]  ( .D(n2738), .CP(clk), .Q(\mem[120][5] ) );
  DFQD1 \mem_reg[120][4]  ( .D(n2737), .CP(clk), .Q(\mem[120][4] ) );
  DFQD1 \mem_reg[120][3]  ( .D(n2736), .CP(clk), .Q(\mem[120][3] ) );
  DFQD1 \mem_reg[120][2]  ( .D(n2735), .CP(clk), .Q(\mem[120][2] ) );
  DFQD1 \mem_reg[120][1]  ( .D(n2734), .CP(clk), .Q(\mem[120][1] ) );
  DFQD1 \mem_reg[120][0]  ( .D(n2733), .CP(clk), .Q(\mem[120][0] ) );
  DFQD1 \mem_reg[121][15]  ( .D(n2732), .CP(clk), .Q(\mem[121][15] ) );
  DFQD1 \mem_reg[121][14]  ( .D(n2731), .CP(clk), .Q(\mem[121][14] ) );
  DFQD1 \mem_reg[121][13]  ( .D(n2730), .CP(clk), .Q(\mem[121][13] ) );
  DFQD1 \mem_reg[121][12]  ( .D(n2729), .CP(clk), .Q(\mem[121][12] ) );
  DFQD1 \mem_reg[121][11]  ( .D(n2728), .CP(clk), .Q(\mem[121][11] ) );
  DFQD1 \mem_reg[121][10]  ( .D(n2727), .CP(clk), .Q(\mem[121][10] ) );
  DFQD1 \mem_reg[121][9]  ( .D(n2726), .CP(clk), .Q(\mem[121][9] ) );
  DFQD1 \mem_reg[121][8]  ( .D(n2725), .CP(clk), .Q(\mem[121][8] ) );
  DFQD1 \mem_reg[121][7]  ( .D(n2724), .CP(clk), .Q(\mem[121][7] ) );
  DFQD1 \mem_reg[121][6]  ( .D(n2723), .CP(clk), .Q(\mem[121][6] ) );
  DFQD1 \mem_reg[121][5]  ( .D(n2722), .CP(clk), .Q(\mem[121][5] ) );
  DFQD1 \mem_reg[121][4]  ( .D(n2721), .CP(clk), .Q(\mem[121][4] ) );
  DFQD1 \mem_reg[121][3]  ( .D(n2720), .CP(clk), .Q(\mem[121][3] ) );
  DFQD1 \mem_reg[121][2]  ( .D(n2719), .CP(clk), .Q(\mem[121][2] ) );
  DFQD1 \mem_reg[121][1]  ( .D(n2718), .CP(clk), .Q(\mem[121][1] ) );
  DFQD1 \mem_reg[121][0]  ( .D(n2717), .CP(clk), .Q(\mem[121][0] ) );
  DFQD1 \mem_reg[122][15]  ( .D(n2716), .CP(clk), .Q(\mem[122][15] ) );
  DFQD1 \mem_reg[122][14]  ( .D(n2715), .CP(clk), .Q(\mem[122][14] ) );
  DFQD1 \mem_reg[122][13]  ( .D(n2714), .CP(clk), .Q(\mem[122][13] ) );
  DFQD1 \mem_reg[122][12]  ( .D(n2713), .CP(clk), .Q(\mem[122][12] ) );
  DFQD1 \mem_reg[122][11]  ( .D(n2712), .CP(clk), .Q(\mem[122][11] ) );
  DFQD1 \mem_reg[122][10]  ( .D(n2711), .CP(clk), .Q(\mem[122][10] ) );
  DFQD1 \mem_reg[122][9]  ( .D(n2710), .CP(clk), .Q(\mem[122][9] ) );
  DFQD1 \mem_reg[122][8]  ( .D(n2709), .CP(clk), .Q(\mem[122][8] ) );
  DFQD1 \mem_reg[122][7]  ( .D(n2708), .CP(clk), .Q(\mem[122][7] ) );
  DFQD1 \mem_reg[122][6]  ( .D(n2707), .CP(clk), .Q(\mem[122][6] ) );
  DFQD1 \mem_reg[122][5]  ( .D(n2706), .CP(clk), .Q(\mem[122][5] ) );
  DFQD1 \mem_reg[122][4]  ( .D(n2705), .CP(clk), .Q(\mem[122][4] ) );
  DFQD1 \mem_reg[122][3]  ( .D(n2704), .CP(clk), .Q(\mem[122][3] ) );
  DFQD1 \mem_reg[122][2]  ( .D(n2703), .CP(clk), .Q(\mem[122][2] ) );
  DFQD1 \mem_reg[122][1]  ( .D(n2702), .CP(clk), .Q(\mem[122][1] ) );
  DFQD1 \mem_reg[122][0]  ( .D(n2701), .CP(clk), .Q(\mem[122][0] ) );
  DFQD1 \mem_reg[123][15]  ( .D(n2700), .CP(clk), .Q(\mem[123][15] ) );
  DFQD1 \mem_reg[123][14]  ( .D(n2699), .CP(clk), .Q(\mem[123][14] ) );
  DFQD1 \mem_reg[123][13]  ( .D(n2698), .CP(clk), .Q(\mem[123][13] ) );
  DFQD1 \mem_reg[123][12]  ( .D(n2697), .CP(clk), .Q(\mem[123][12] ) );
  DFQD1 \mem_reg[123][11]  ( .D(n2696), .CP(clk), .Q(\mem[123][11] ) );
  DFQD1 \mem_reg[123][10]  ( .D(n2695), .CP(clk), .Q(\mem[123][10] ) );
  DFQD1 \mem_reg[123][9]  ( .D(n2694), .CP(clk), .Q(\mem[123][9] ) );
  DFQD1 \mem_reg[123][8]  ( .D(n2693), .CP(clk), .Q(\mem[123][8] ) );
  DFQD1 \mem_reg[123][7]  ( .D(n2692), .CP(clk), .Q(\mem[123][7] ) );
  DFQD1 \mem_reg[123][6]  ( .D(n2691), .CP(clk), .Q(\mem[123][6] ) );
  DFQD1 \mem_reg[123][5]  ( .D(n2690), .CP(clk), .Q(\mem[123][5] ) );
  DFQD1 \mem_reg[123][4]  ( .D(n2689), .CP(clk), .Q(\mem[123][4] ) );
  DFQD1 \mem_reg[123][3]  ( .D(n2688), .CP(clk), .Q(\mem[123][3] ) );
  DFQD1 \mem_reg[123][2]  ( .D(n2687), .CP(clk), .Q(\mem[123][2] ) );
  DFQD1 \mem_reg[123][1]  ( .D(n2686), .CP(clk), .Q(\mem[123][1] ) );
  DFQD1 \mem_reg[123][0]  ( .D(n2685), .CP(clk), .Q(\mem[123][0] ) );
  DFQD1 \mem_reg[124][15]  ( .D(n2684), .CP(clk), .Q(\mem[124][15] ) );
  DFQD1 \mem_reg[124][14]  ( .D(n2683), .CP(clk), .Q(\mem[124][14] ) );
  DFQD1 \mem_reg[124][13]  ( .D(n2682), .CP(clk), .Q(\mem[124][13] ) );
  DFQD1 \mem_reg[124][12]  ( .D(n2681), .CP(clk), .Q(\mem[124][12] ) );
  DFQD1 \mem_reg[124][11]  ( .D(n2680), .CP(clk), .Q(\mem[124][11] ) );
  DFQD1 \mem_reg[124][10]  ( .D(n2679), .CP(clk), .Q(\mem[124][10] ) );
  DFQD1 \mem_reg[124][9]  ( .D(n2678), .CP(clk), .Q(\mem[124][9] ) );
  DFQD1 \mem_reg[124][8]  ( .D(n2677), .CP(clk), .Q(\mem[124][8] ) );
  DFQD1 \mem_reg[124][7]  ( .D(n2676), .CP(clk), .Q(\mem[124][7] ) );
  DFQD1 \mem_reg[124][6]  ( .D(n2675), .CP(clk), .Q(\mem[124][6] ) );
  DFQD1 \mem_reg[124][5]  ( .D(n2674), .CP(clk), .Q(\mem[124][5] ) );
  DFQD1 \mem_reg[124][4]  ( .D(n2673), .CP(clk), .Q(\mem[124][4] ) );
  DFQD1 \mem_reg[124][3]  ( .D(n2672), .CP(clk), .Q(\mem[124][3] ) );
  DFQD1 \mem_reg[124][2]  ( .D(n2671), .CP(clk), .Q(\mem[124][2] ) );
  DFQD1 \mem_reg[124][1]  ( .D(n2670), .CP(clk), .Q(\mem[124][1] ) );
  DFQD1 \mem_reg[124][0]  ( .D(n2669), .CP(clk), .Q(\mem[124][0] ) );
  DFQD1 \mem_reg[125][15]  ( .D(n2668), .CP(clk), .Q(\mem[125][15] ) );
  DFQD1 \mem_reg[125][14]  ( .D(n2667), .CP(clk), .Q(\mem[125][14] ) );
  DFQD1 \mem_reg[125][13]  ( .D(n2666), .CP(clk), .Q(\mem[125][13] ) );
  DFQD1 \mem_reg[125][12]  ( .D(n2665), .CP(clk), .Q(\mem[125][12] ) );
  DFQD1 \mem_reg[125][11]  ( .D(n2664), .CP(clk), .Q(\mem[125][11] ) );
  DFQD1 \mem_reg[125][10]  ( .D(n2663), .CP(clk), .Q(\mem[125][10] ) );
  DFQD1 \mem_reg[125][9]  ( .D(n2662), .CP(clk), .Q(\mem[125][9] ) );
  DFQD1 \mem_reg[125][8]  ( .D(n2661), .CP(clk), .Q(\mem[125][8] ) );
  DFQD1 \mem_reg[125][7]  ( .D(n2660), .CP(clk), .Q(\mem[125][7] ) );
  DFQD1 \mem_reg[125][6]  ( .D(n2659), .CP(clk), .Q(\mem[125][6] ) );
  DFQD1 \mem_reg[125][5]  ( .D(n2658), .CP(clk), .Q(\mem[125][5] ) );
  DFQD1 \mem_reg[125][4]  ( .D(n2657), .CP(clk), .Q(\mem[125][4] ) );
  DFQD1 \mem_reg[125][3]  ( .D(n2656), .CP(clk), .Q(\mem[125][3] ) );
  DFQD1 \mem_reg[125][2]  ( .D(n2655), .CP(clk), .Q(\mem[125][2] ) );
  DFQD1 \mem_reg[125][1]  ( .D(n2654), .CP(clk), .Q(\mem[125][1] ) );
  DFQD1 \mem_reg[125][0]  ( .D(n2653), .CP(clk), .Q(\mem[125][0] ) );
  DFQD1 \mem_reg[126][15]  ( .D(n2652), .CP(clk), .Q(\mem[126][15] ) );
  DFQD1 \mem_reg[126][14]  ( .D(n2651), .CP(clk), .Q(\mem[126][14] ) );
  DFQD1 \mem_reg[126][13]  ( .D(n2650), .CP(clk), .Q(\mem[126][13] ) );
  DFQD1 \mem_reg[126][12]  ( .D(n2649), .CP(clk), .Q(\mem[126][12] ) );
  DFQD1 \mem_reg[126][11]  ( .D(n2648), .CP(clk), .Q(\mem[126][11] ) );
  DFQD1 \mem_reg[126][10]  ( .D(n2647), .CP(clk), .Q(\mem[126][10] ) );
  DFQD1 \mem_reg[126][9]  ( .D(n2646), .CP(clk), .Q(\mem[126][9] ) );
  DFQD1 \mem_reg[126][8]  ( .D(n2645), .CP(clk), .Q(\mem[126][8] ) );
  DFQD1 \mem_reg[126][7]  ( .D(n2644), .CP(clk), .Q(\mem[126][7] ) );
  DFQD1 \mem_reg[126][6]  ( .D(n2643), .CP(clk), .Q(\mem[126][6] ) );
  DFQD1 \mem_reg[126][5]  ( .D(n2642), .CP(clk), .Q(\mem[126][5] ) );
  DFQD1 \mem_reg[126][4]  ( .D(n2641), .CP(clk), .Q(\mem[126][4] ) );
  DFQD1 \mem_reg[126][3]  ( .D(n2640), .CP(clk), .Q(\mem[126][3] ) );
  DFQD1 \mem_reg[126][2]  ( .D(n2639), .CP(clk), .Q(\mem[126][2] ) );
  DFQD1 \mem_reg[126][1]  ( .D(n2638), .CP(clk), .Q(\mem[126][1] ) );
  DFQD1 \mem_reg[126][0]  ( .D(n2637), .CP(clk), .Q(\mem[126][0] ) );
  DFQD1 \mem_reg[127][15]  ( .D(n2636), .CP(clk), .Q(\mem[127][15] ) );
  DFQD1 \mem_reg[127][14]  ( .D(n2635), .CP(clk), .Q(\mem[127][14] ) );
  DFQD1 \mem_reg[127][13]  ( .D(n2634), .CP(clk), .Q(\mem[127][13] ) );
  DFQD1 \mem_reg[127][12]  ( .D(n2633), .CP(clk), .Q(\mem[127][12] ) );
  DFQD1 \mem_reg[127][11]  ( .D(n2632), .CP(clk), .Q(\mem[127][11] ) );
  DFQD1 \mem_reg[127][10]  ( .D(n2631), .CP(clk), .Q(\mem[127][10] ) );
  DFQD1 \mem_reg[127][9]  ( .D(n2630), .CP(clk), .Q(\mem[127][9] ) );
  DFQD1 \mem_reg[127][8]  ( .D(n2629), .CP(clk), .Q(\mem[127][8] ) );
  DFQD1 \mem_reg[127][7]  ( .D(n2628), .CP(clk), .Q(\mem[127][7] ) );
  DFQD1 \mem_reg[127][6]  ( .D(n2627), .CP(clk), .Q(\mem[127][6] ) );
  DFQD1 \mem_reg[127][5]  ( .D(n2626), .CP(clk), .Q(\mem[127][5] ) );
  DFQD1 \mem_reg[127][4]  ( .D(n2625), .CP(clk), .Q(\mem[127][4] ) );
  DFQD1 \mem_reg[127][3]  ( .D(n2624), .CP(clk), .Q(\mem[127][3] ) );
  DFQD1 \mem_reg[127][2]  ( .D(n2623), .CP(clk), .Q(\mem[127][2] ) );
  DFQD1 \mem_reg[127][1]  ( .D(n2622), .CP(clk), .Q(\mem[127][1] ) );
  DFQD1 \mem_reg[127][0]  ( .D(n2621), .CP(clk), .Q(\mem[127][0] ) );
  DFQD1 \mem_reg[128][15]  ( .D(n2620), .CP(clk), .Q(\mem[128][15] ) );
  DFQD1 \mem_reg[128][14]  ( .D(n2619), .CP(clk), .Q(\mem[128][14] ) );
  DFQD1 \mem_reg[128][13]  ( .D(n2618), .CP(clk), .Q(\mem[128][13] ) );
  DFQD1 \mem_reg[128][12]  ( .D(n2617), .CP(clk), .Q(\mem[128][12] ) );
  DFQD1 \mem_reg[128][11]  ( .D(n2616), .CP(clk), .Q(\mem[128][11] ) );
  DFQD1 \mem_reg[128][10]  ( .D(n2615), .CP(clk), .Q(\mem[128][10] ) );
  DFQD1 \mem_reg[128][9]  ( .D(n2614), .CP(clk), .Q(\mem[128][9] ) );
  DFQD1 \mem_reg[128][8]  ( .D(n2613), .CP(clk), .Q(\mem[128][8] ) );
  DFQD1 \mem_reg[128][7]  ( .D(n2612), .CP(clk), .Q(\mem[128][7] ) );
  DFQD1 \mem_reg[128][6]  ( .D(n2611), .CP(clk), .Q(\mem[128][6] ) );
  DFQD1 \mem_reg[128][5]  ( .D(n2610), .CP(clk), .Q(\mem[128][5] ) );
  DFQD1 \mem_reg[128][4]  ( .D(n2609), .CP(clk), .Q(\mem[128][4] ) );
  DFQD1 \mem_reg[128][3]  ( .D(n2608), .CP(clk), .Q(\mem[128][3] ) );
  DFQD1 \mem_reg[128][2]  ( .D(n2607), .CP(clk), .Q(\mem[128][2] ) );
  DFQD1 \mem_reg[128][1]  ( .D(n2606), .CP(clk), .Q(\mem[128][1] ) );
  DFQD1 \mem_reg[128][0]  ( .D(n2605), .CP(clk), .Q(\mem[128][0] ) );
  DFQD1 \mem_reg[129][15]  ( .D(n2604), .CP(clk), .Q(\mem[129][15] ) );
  DFQD1 \mem_reg[129][14]  ( .D(n2603), .CP(clk), .Q(\mem[129][14] ) );
  DFQD1 \mem_reg[129][13]  ( .D(n2602), .CP(clk), .Q(\mem[129][13] ) );
  DFQD1 \mem_reg[129][12]  ( .D(n2601), .CP(clk), .Q(\mem[129][12] ) );
  DFQD1 \mem_reg[129][11]  ( .D(n2600), .CP(clk), .Q(\mem[129][11] ) );
  DFQD1 \mem_reg[129][10]  ( .D(n2599), .CP(clk), .Q(\mem[129][10] ) );
  DFQD1 \mem_reg[129][9]  ( .D(n2598), .CP(clk), .Q(\mem[129][9] ) );
  DFQD1 \mem_reg[129][8]  ( .D(n2597), .CP(clk), .Q(\mem[129][8] ) );
  DFQD1 \mem_reg[129][7]  ( .D(n2596), .CP(clk), .Q(\mem[129][7] ) );
  DFQD1 \mem_reg[129][6]  ( .D(n2595), .CP(clk), .Q(\mem[129][6] ) );
  DFQD1 \mem_reg[129][5]  ( .D(n2594), .CP(clk), .Q(\mem[129][5] ) );
  DFQD1 \mem_reg[129][4]  ( .D(n2593), .CP(clk), .Q(\mem[129][4] ) );
  DFQD1 \mem_reg[129][3]  ( .D(n2592), .CP(clk), .Q(\mem[129][3] ) );
  DFQD1 \mem_reg[129][2]  ( .D(n2591), .CP(clk), .Q(\mem[129][2] ) );
  DFQD1 \mem_reg[129][1]  ( .D(n2590), .CP(clk), .Q(\mem[129][1] ) );
  DFQD1 \mem_reg[129][0]  ( .D(n2589), .CP(clk), .Q(\mem[129][0] ) );
  DFQD1 \mem_reg[130][15]  ( .D(n2588), .CP(clk), .Q(\mem[130][15] ) );
  DFQD1 \mem_reg[130][14]  ( .D(n2587), .CP(clk), .Q(\mem[130][14] ) );
  DFQD1 \mem_reg[130][13]  ( .D(n2586), .CP(clk), .Q(\mem[130][13] ) );
  DFQD1 \mem_reg[130][12]  ( .D(n2585), .CP(clk), .Q(\mem[130][12] ) );
  DFQD1 \mem_reg[130][11]  ( .D(n2584), .CP(clk), .Q(\mem[130][11] ) );
  DFQD1 \mem_reg[130][10]  ( .D(n2583), .CP(clk), .Q(\mem[130][10] ) );
  DFQD1 \mem_reg[130][9]  ( .D(n2582), .CP(clk), .Q(\mem[130][9] ) );
  DFQD1 \mem_reg[130][8]  ( .D(n2581), .CP(clk), .Q(\mem[130][8] ) );
  DFQD1 \mem_reg[130][7]  ( .D(n2580), .CP(clk), .Q(\mem[130][7] ) );
  DFQD1 \mem_reg[130][6]  ( .D(n2579), .CP(clk), .Q(\mem[130][6] ) );
  DFQD1 \mem_reg[130][5]  ( .D(n2578), .CP(clk), .Q(\mem[130][5] ) );
  DFQD1 \mem_reg[130][4]  ( .D(n2577), .CP(clk), .Q(\mem[130][4] ) );
  DFQD1 \mem_reg[130][3]  ( .D(n2576), .CP(clk), .Q(\mem[130][3] ) );
  DFQD1 \mem_reg[130][2]  ( .D(n2575), .CP(clk), .Q(\mem[130][2] ) );
  DFQD1 \mem_reg[130][1]  ( .D(n2574), .CP(clk), .Q(\mem[130][1] ) );
  DFQD1 \mem_reg[130][0]  ( .D(n2573), .CP(clk), .Q(\mem[130][0] ) );
  DFQD1 \mem_reg[131][15]  ( .D(n2572), .CP(clk), .Q(\mem[131][15] ) );
  DFQD1 \mem_reg[131][14]  ( .D(n2571), .CP(clk), .Q(\mem[131][14] ) );
  DFQD1 \mem_reg[131][13]  ( .D(n2570), .CP(clk), .Q(\mem[131][13] ) );
  DFQD1 \mem_reg[131][12]  ( .D(n2569), .CP(clk), .Q(\mem[131][12] ) );
  DFQD1 \mem_reg[131][11]  ( .D(n2568), .CP(clk), .Q(\mem[131][11] ) );
  DFQD1 \mem_reg[131][10]  ( .D(n2567), .CP(clk), .Q(\mem[131][10] ) );
  DFQD1 \mem_reg[131][9]  ( .D(n2566), .CP(clk), .Q(\mem[131][9] ) );
  DFQD1 \mem_reg[131][8]  ( .D(n2565), .CP(clk), .Q(\mem[131][8] ) );
  DFQD1 \mem_reg[131][7]  ( .D(n2564), .CP(clk), .Q(\mem[131][7] ) );
  DFQD1 \mem_reg[131][6]  ( .D(n2563), .CP(clk), .Q(\mem[131][6] ) );
  DFQD1 \mem_reg[131][5]  ( .D(n2562), .CP(clk), .Q(\mem[131][5] ) );
  DFQD1 \mem_reg[131][4]  ( .D(n2561), .CP(clk), .Q(\mem[131][4] ) );
  DFQD1 \mem_reg[131][3]  ( .D(n2560), .CP(clk), .Q(\mem[131][3] ) );
  DFQD1 \mem_reg[131][2]  ( .D(n2559), .CP(clk), .Q(\mem[131][2] ) );
  DFQD1 \mem_reg[131][1]  ( .D(n2558), .CP(clk), .Q(\mem[131][1] ) );
  DFQD1 \mem_reg[131][0]  ( .D(n2557), .CP(clk), .Q(\mem[131][0] ) );
  DFQD1 \mem_reg[132][15]  ( .D(n2556), .CP(clk), .Q(\mem[132][15] ) );
  DFQD1 \mem_reg[132][14]  ( .D(n2555), .CP(clk), .Q(\mem[132][14] ) );
  DFQD1 \mem_reg[132][13]  ( .D(n2554), .CP(clk), .Q(\mem[132][13] ) );
  DFQD1 \mem_reg[132][12]  ( .D(n2553), .CP(clk), .Q(\mem[132][12] ) );
  DFQD1 \mem_reg[132][11]  ( .D(n2552), .CP(clk), .Q(\mem[132][11] ) );
  DFQD1 \mem_reg[132][10]  ( .D(n2551), .CP(clk), .Q(\mem[132][10] ) );
  DFQD1 \mem_reg[132][9]  ( .D(n2550), .CP(clk), .Q(\mem[132][9] ) );
  DFQD1 \mem_reg[132][8]  ( .D(n2549), .CP(clk), .Q(\mem[132][8] ) );
  DFQD1 \mem_reg[132][7]  ( .D(n2548), .CP(clk), .Q(\mem[132][7] ) );
  DFQD1 \mem_reg[132][6]  ( .D(n2547), .CP(clk), .Q(\mem[132][6] ) );
  DFQD1 \mem_reg[132][5]  ( .D(n2546), .CP(clk), .Q(\mem[132][5] ) );
  DFQD1 \mem_reg[132][4]  ( .D(n2545), .CP(clk), .Q(\mem[132][4] ) );
  DFQD1 \mem_reg[132][3]  ( .D(n2544), .CP(clk), .Q(\mem[132][3] ) );
  DFQD1 \mem_reg[132][2]  ( .D(n2543), .CP(clk), .Q(\mem[132][2] ) );
  DFQD1 \mem_reg[132][1]  ( .D(n2542), .CP(clk), .Q(\mem[132][1] ) );
  DFQD1 \mem_reg[132][0]  ( .D(n2541), .CP(clk), .Q(\mem[132][0] ) );
  DFQD1 \mem_reg[133][15]  ( .D(n2540), .CP(clk), .Q(\mem[133][15] ) );
  DFQD1 \mem_reg[133][14]  ( .D(n2539), .CP(clk), .Q(\mem[133][14] ) );
  DFQD1 \mem_reg[133][13]  ( .D(n2538), .CP(clk), .Q(\mem[133][13] ) );
  DFQD1 \mem_reg[133][12]  ( .D(n2537), .CP(clk), .Q(\mem[133][12] ) );
  DFQD1 \mem_reg[133][11]  ( .D(n2536), .CP(clk), .Q(\mem[133][11] ) );
  DFQD1 \mem_reg[133][10]  ( .D(n2535), .CP(clk), .Q(\mem[133][10] ) );
  DFQD1 \mem_reg[133][9]  ( .D(n2534), .CP(clk), .Q(\mem[133][9] ) );
  DFQD1 \mem_reg[133][8]  ( .D(n2533), .CP(clk), .Q(\mem[133][8] ) );
  DFQD1 \mem_reg[133][7]  ( .D(n2532), .CP(clk), .Q(\mem[133][7] ) );
  DFQD1 \mem_reg[133][6]  ( .D(n2531), .CP(clk), .Q(\mem[133][6] ) );
  DFQD1 \mem_reg[133][5]  ( .D(n2530), .CP(clk), .Q(\mem[133][5] ) );
  DFQD1 \mem_reg[133][4]  ( .D(n2529), .CP(clk), .Q(\mem[133][4] ) );
  DFQD1 \mem_reg[133][3]  ( .D(n2528), .CP(clk), .Q(\mem[133][3] ) );
  DFQD1 \mem_reg[133][2]  ( .D(n2527), .CP(clk), .Q(\mem[133][2] ) );
  DFQD1 \mem_reg[133][1]  ( .D(n2526), .CP(clk), .Q(\mem[133][1] ) );
  DFQD1 \mem_reg[133][0]  ( .D(n2525), .CP(clk), .Q(\mem[133][0] ) );
  DFQD1 \mem_reg[134][15]  ( .D(n2524), .CP(clk), .Q(\mem[134][15] ) );
  DFQD1 \mem_reg[134][14]  ( .D(n2523), .CP(clk), .Q(\mem[134][14] ) );
  DFQD1 \mem_reg[134][13]  ( .D(n2522), .CP(clk), .Q(\mem[134][13] ) );
  DFQD1 \mem_reg[134][12]  ( .D(n2521), .CP(clk), .Q(\mem[134][12] ) );
  DFQD1 \mem_reg[134][11]  ( .D(n2520), .CP(clk), .Q(\mem[134][11] ) );
  DFQD1 \mem_reg[134][10]  ( .D(n2519), .CP(clk), .Q(\mem[134][10] ) );
  DFQD1 \mem_reg[134][9]  ( .D(n2518), .CP(clk), .Q(\mem[134][9] ) );
  DFQD1 \mem_reg[134][8]  ( .D(n2517), .CP(clk), .Q(\mem[134][8] ) );
  DFQD1 \mem_reg[134][7]  ( .D(n2516), .CP(clk), .Q(\mem[134][7] ) );
  DFQD1 \mem_reg[134][6]  ( .D(n2515), .CP(clk), .Q(\mem[134][6] ) );
  DFQD1 \mem_reg[134][5]  ( .D(n2514), .CP(clk), .Q(\mem[134][5] ) );
  DFQD1 \mem_reg[134][4]  ( .D(n2513), .CP(clk), .Q(\mem[134][4] ) );
  DFQD1 \mem_reg[134][3]  ( .D(n2512), .CP(clk), .Q(\mem[134][3] ) );
  DFQD1 \mem_reg[134][2]  ( .D(n2511), .CP(clk), .Q(\mem[134][2] ) );
  DFQD1 \mem_reg[134][1]  ( .D(n2510), .CP(clk), .Q(\mem[134][1] ) );
  DFQD1 \mem_reg[134][0]  ( .D(n2509), .CP(clk), .Q(\mem[134][0] ) );
  DFQD1 \mem_reg[135][15]  ( .D(n2508), .CP(clk), .Q(\mem[135][15] ) );
  DFQD1 \mem_reg[135][14]  ( .D(n2507), .CP(clk), .Q(\mem[135][14] ) );
  DFQD1 \mem_reg[135][13]  ( .D(n2506), .CP(clk), .Q(\mem[135][13] ) );
  DFQD1 \mem_reg[135][12]  ( .D(n2505), .CP(clk), .Q(\mem[135][12] ) );
  DFQD1 \mem_reg[135][11]  ( .D(n2504), .CP(clk), .Q(\mem[135][11] ) );
  DFQD1 \mem_reg[135][10]  ( .D(n2503), .CP(clk), .Q(\mem[135][10] ) );
  DFQD1 \mem_reg[135][9]  ( .D(n2502), .CP(clk), .Q(\mem[135][9] ) );
  DFQD1 \mem_reg[135][8]  ( .D(n2501), .CP(clk), .Q(\mem[135][8] ) );
  DFQD1 \mem_reg[135][7]  ( .D(n2500), .CP(clk), .Q(\mem[135][7] ) );
  DFQD1 \mem_reg[135][6]  ( .D(n2499), .CP(clk), .Q(\mem[135][6] ) );
  DFQD1 \mem_reg[135][5]  ( .D(n2498), .CP(clk), .Q(\mem[135][5] ) );
  DFQD1 \mem_reg[135][4]  ( .D(n2497), .CP(clk), .Q(\mem[135][4] ) );
  DFQD1 \mem_reg[135][3]  ( .D(n2496), .CP(clk), .Q(\mem[135][3] ) );
  DFQD1 \mem_reg[135][2]  ( .D(n2495), .CP(clk), .Q(\mem[135][2] ) );
  DFQD1 \mem_reg[135][1]  ( .D(n2494), .CP(clk), .Q(\mem[135][1] ) );
  DFQD1 \mem_reg[135][0]  ( .D(n2493), .CP(clk), .Q(\mem[135][0] ) );
  DFQD1 \mem_reg[136][15]  ( .D(n2492), .CP(clk), .Q(\mem[136][15] ) );
  DFQD1 \mem_reg[136][14]  ( .D(n2491), .CP(clk), .Q(\mem[136][14] ) );
  DFQD1 \mem_reg[136][13]  ( .D(n2490), .CP(clk), .Q(\mem[136][13] ) );
  DFQD1 \mem_reg[136][12]  ( .D(n2489), .CP(clk), .Q(\mem[136][12] ) );
  DFQD1 \mem_reg[136][11]  ( .D(n2488), .CP(clk), .Q(\mem[136][11] ) );
  DFQD1 \mem_reg[136][10]  ( .D(n2487), .CP(clk), .Q(\mem[136][10] ) );
  DFQD1 \mem_reg[136][9]  ( .D(n2486), .CP(clk), .Q(\mem[136][9] ) );
  DFQD1 \mem_reg[136][8]  ( .D(n2485), .CP(clk), .Q(\mem[136][8] ) );
  DFQD1 \mem_reg[136][7]  ( .D(n2484), .CP(clk), .Q(\mem[136][7] ) );
  DFQD1 \mem_reg[136][6]  ( .D(n2483), .CP(clk), .Q(\mem[136][6] ) );
  DFQD1 \mem_reg[136][5]  ( .D(n2482), .CP(clk), .Q(\mem[136][5] ) );
  DFQD1 \mem_reg[136][4]  ( .D(n2481), .CP(clk), .Q(\mem[136][4] ) );
  DFQD1 \mem_reg[136][3]  ( .D(n2480), .CP(clk), .Q(\mem[136][3] ) );
  DFQD1 \mem_reg[136][2]  ( .D(n2479), .CP(clk), .Q(\mem[136][2] ) );
  DFQD1 \mem_reg[136][1]  ( .D(n2478), .CP(clk), .Q(\mem[136][1] ) );
  DFQD1 \mem_reg[136][0]  ( .D(n2477), .CP(clk), .Q(\mem[136][0] ) );
  DFQD1 \mem_reg[137][15]  ( .D(n2476), .CP(clk), .Q(\mem[137][15] ) );
  DFQD1 \mem_reg[137][14]  ( .D(n2475), .CP(clk), .Q(\mem[137][14] ) );
  DFQD1 \mem_reg[137][13]  ( .D(n2474), .CP(clk), .Q(\mem[137][13] ) );
  DFQD1 \mem_reg[137][12]  ( .D(n2473), .CP(clk), .Q(\mem[137][12] ) );
  DFQD1 \mem_reg[137][11]  ( .D(n2472), .CP(clk), .Q(\mem[137][11] ) );
  DFQD1 \mem_reg[137][10]  ( .D(n2471), .CP(clk), .Q(\mem[137][10] ) );
  DFQD1 \mem_reg[137][9]  ( .D(n2470), .CP(clk), .Q(\mem[137][9] ) );
  DFQD1 \mem_reg[137][8]  ( .D(n2469), .CP(clk), .Q(\mem[137][8] ) );
  DFQD1 \mem_reg[137][7]  ( .D(n2468), .CP(clk), .Q(\mem[137][7] ) );
  DFQD1 \mem_reg[137][6]  ( .D(n2467), .CP(clk), .Q(\mem[137][6] ) );
  DFQD1 \mem_reg[137][5]  ( .D(n2466), .CP(clk), .Q(\mem[137][5] ) );
  DFQD1 \mem_reg[137][4]  ( .D(n2465), .CP(clk), .Q(\mem[137][4] ) );
  DFQD1 \mem_reg[137][3]  ( .D(n2464), .CP(clk), .Q(\mem[137][3] ) );
  DFQD1 \mem_reg[137][2]  ( .D(n2463), .CP(clk), .Q(\mem[137][2] ) );
  DFQD1 \mem_reg[137][1]  ( .D(n2462), .CP(clk), .Q(\mem[137][1] ) );
  DFQD1 \mem_reg[137][0]  ( .D(n2461), .CP(clk), .Q(\mem[137][0] ) );
  DFQD1 \mem_reg[138][15]  ( .D(n2460), .CP(clk), .Q(\mem[138][15] ) );
  DFQD1 \mem_reg[138][14]  ( .D(n2459), .CP(clk), .Q(\mem[138][14] ) );
  DFQD1 \mem_reg[138][13]  ( .D(n2458), .CP(clk), .Q(\mem[138][13] ) );
  DFQD1 \mem_reg[138][12]  ( .D(n2457), .CP(clk), .Q(\mem[138][12] ) );
  DFQD1 \mem_reg[138][11]  ( .D(n2456), .CP(clk), .Q(\mem[138][11] ) );
  DFQD1 \mem_reg[138][10]  ( .D(n2455), .CP(clk), .Q(\mem[138][10] ) );
  DFQD1 \mem_reg[138][9]  ( .D(n2454), .CP(clk), .Q(\mem[138][9] ) );
  DFQD1 \mem_reg[138][8]  ( .D(n2453), .CP(clk), .Q(\mem[138][8] ) );
  DFQD1 \mem_reg[138][7]  ( .D(n2452), .CP(clk), .Q(\mem[138][7] ) );
  DFQD1 \mem_reg[138][6]  ( .D(n2451), .CP(clk), .Q(\mem[138][6] ) );
  DFQD1 \mem_reg[138][5]  ( .D(n2450), .CP(clk), .Q(\mem[138][5] ) );
  DFQD1 \mem_reg[138][4]  ( .D(n2449), .CP(clk), .Q(\mem[138][4] ) );
  DFQD1 \mem_reg[138][3]  ( .D(n2448), .CP(clk), .Q(\mem[138][3] ) );
  DFQD1 \mem_reg[138][2]  ( .D(n2447), .CP(clk), .Q(\mem[138][2] ) );
  DFQD1 \mem_reg[138][1]  ( .D(n2446), .CP(clk), .Q(\mem[138][1] ) );
  DFQD1 \mem_reg[138][0]  ( .D(n2445), .CP(clk), .Q(\mem[138][0] ) );
  DFQD1 \mem_reg[139][15]  ( .D(n2444), .CP(clk), .Q(\mem[139][15] ) );
  DFQD1 \mem_reg[139][14]  ( .D(n2443), .CP(clk), .Q(\mem[139][14] ) );
  DFQD1 \mem_reg[139][13]  ( .D(n2442), .CP(clk), .Q(\mem[139][13] ) );
  DFQD1 \mem_reg[139][12]  ( .D(n2441), .CP(clk), .Q(\mem[139][12] ) );
  DFQD1 \mem_reg[139][11]  ( .D(n2440), .CP(clk), .Q(\mem[139][11] ) );
  DFQD1 \mem_reg[139][10]  ( .D(n2439), .CP(clk), .Q(\mem[139][10] ) );
  DFQD1 \mem_reg[139][9]  ( .D(n2438), .CP(clk), .Q(\mem[139][9] ) );
  DFQD1 \mem_reg[139][8]  ( .D(n2437), .CP(clk), .Q(\mem[139][8] ) );
  DFQD1 \mem_reg[139][7]  ( .D(n2436), .CP(clk), .Q(\mem[139][7] ) );
  DFQD1 \mem_reg[139][6]  ( .D(n2435), .CP(clk), .Q(\mem[139][6] ) );
  DFQD1 \mem_reg[139][5]  ( .D(n2434), .CP(clk), .Q(\mem[139][5] ) );
  DFQD1 \mem_reg[139][4]  ( .D(n2433), .CP(clk), .Q(\mem[139][4] ) );
  DFQD1 \mem_reg[139][3]  ( .D(n2432), .CP(clk), .Q(\mem[139][3] ) );
  DFQD1 \mem_reg[139][2]  ( .D(n2431), .CP(clk), .Q(\mem[139][2] ) );
  DFQD1 \mem_reg[139][1]  ( .D(n2430), .CP(clk), .Q(\mem[139][1] ) );
  DFQD1 \mem_reg[139][0]  ( .D(n2429), .CP(clk), .Q(\mem[139][0] ) );
  DFQD1 \mem_reg[140][15]  ( .D(n2428), .CP(clk), .Q(\mem[140][15] ) );
  DFQD1 \mem_reg[140][14]  ( .D(n2427), .CP(clk), .Q(\mem[140][14] ) );
  DFQD1 \mem_reg[140][13]  ( .D(n2426), .CP(clk), .Q(\mem[140][13] ) );
  DFQD1 \mem_reg[140][12]  ( .D(n2425), .CP(clk), .Q(\mem[140][12] ) );
  DFQD1 \mem_reg[140][11]  ( .D(n2424), .CP(clk), .Q(\mem[140][11] ) );
  DFQD1 \mem_reg[140][10]  ( .D(n2423), .CP(clk), .Q(\mem[140][10] ) );
  DFQD1 \mem_reg[140][9]  ( .D(n2422), .CP(clk), .Q(\mem[140][9] ) );
  DFQD1 \mem_reg[140][8]  ( .D(n2421), .CP(clk), .Q(\mem[140][8] ) );
  DFQD1 \mem_reg[140][7]  ( .D(n2420), .CP(clk), .Q(\mem[140][7] ) );
  DFQD1 \mem_reg[140][6]  ( .D(n2419), .CP(clk), .Q(\mem[140][6] ) );
  DFQD1 \mem_reg[140][5]  ( .D(n2418), .CP(clk), .Q(\mem[140][5] ) );
  DFQD1 \mem_reg[140][4]  ( .D(n2417), .CP(clk), .Q(\mem[140][4] ) );
  DFQD1 \mem_reg[140][3]  ( .D(n2416), .CP(clk), .Q(\mem[140][3] ) );
  DFQD1 \mem_reg[140][2]  ( .D(n2415), .CP(clk), .Q(\mem[140][2] ) );
  DFQD1 \mem_reg[140][1]  ( .D(n2414), .CP(clk), .Q(\mem[140][1] ) );
  DFQD1 \mem_reg[140][0]  ( .D(n2413), .CP(clk), .Q(\mem[140][0] ) );
  DFQD1 \mem_reg[141][15]  ( .D(n2412), .CP(clk), .Q(\mem[141][15] ) );
  DFQD1 \mem_reg[141][14]  ( .D(n2411), .CP(clk), .Q(\mem[141][14] ) );
  DFQD1 \mem_reg[141][13]  ( .D(n2410), .CP(clk), .Q(\mem[141][13] ) );
  DFQD1 \mem_reg[141][12]  ( .D(n2409), .CP(clk), .Q(\mem[141][12] ) );
  DFQD1 \mem_reg[141][11]  ( .D(n2408), .CP(clk), .Q(\mem[141][11] ) );
  DFQD1 \mem_reg[141][10]  ( .D(n2407), .CP(clk), .Q(\mem[141][10] ) );
  DFQD1 \mem_reg[141][9]  ( .D(n2406), .CP(clk), .Q(\mem[141][9] ) );
  DFQD1 \mem_reg[141][8]  ( .D(n2405), .CP(clk), .Q(\mem[141][8] ) );
  DFQD1 \mem_reg[141][7]  ( .D(n2404), .CP(clk), .Q(\mem[141][7] ) );
  DFQD1 \mem_reg[141][6]  ( .D(n2403), .CP(clk), .Q(\mem[141][6] ) );
  DFQD1 \mem_reg[141][5]  ( .D(n2402), .CP(clk), .Q(\mem[141][5] ) );
  DFQD1 \mem_reg[141][4]  ( .D(n2401), .CP(clk), .Q(\mem[141][4] ) );
  DFQD1 \mem_reg[141][3]  ( .D(n2400), .CP(clk), .Q(\mem[141][3] ) );
  DFQD1 \mem_reg[141][2]  ( .D(n2399), .CP(clk), .Q(\mem[141][2] ) );
  DFQD1 \mem_reg[141][1]  ( .D(n2398), .CP(clk), .Q(\mem[141][1] ) );
  DFQD1 \mem_reg[141][0]  ( .D(n2397), .CP(clk), .Q(\mem[141][0] ) );
  DFQD1 \mem_reg[142][15]  ( .D(n2396), .CP(clk), .Q(\mem[142][15] ) );
  DFQD1 \mem_reg[142][14]  ( .D(n2395), .CP(clk), .Q(\mem[142][14] ) );
  DFQD1 \mem_reg[142][13]  ( .D(n2394), .CP(clk), .Q(\mem[142][13] ) );
  DFQD1 \mem_reg[142][12]  ( .D(n2393), .CP(clk), .Q(\mem[142][12] ) );
  DFQD1 \mem_reg[142][11]  ( .D(n2392), .CP(clk), .Q(\mem[142][11] ) );
  DFQD1 \mem_reg[142][10]  ( .D(n2391), .CP(clk), .Q(\mem[142][10] ) );
  DFQD1 \mem_reg[142][9]  ( .D(n2390), .CP(clk), .Q(\mem[142][9] ) );
  DFQD1 \mem_reg[142][8]  ( .D(n2389), .CP(clk), .Q(\mem[142][8] ) );
  DFQD1 \mem_reg[142][7]  ( .D(n2388), .CP(clk), .Q(\mem[142][7] ) );
  DFQD1 \mem_reg[142][6]  ( .D(n2387), .CP(clk), .Q(\mem[142][6] ) );
  DFQD1 \mem_reg[142][5]  ( .D(n2386), .CP(clk), .Q(\mem[142][5] ) );
  DFQD1 \mem_reg[142][4]  ( .D(n2385), .CP(clk), .Q(\mem[142][4] ) );
  DFQD1 \mem_reg[142][3]  ( .D(n2384), .CP(clk), .Q(\mem[142][3] ) );
  DFQD1 \mem_reg[142][2]  ( .D(n2383), .CP(clk), .Q(\mem[142][2] ) );
  DFQD1 \mem_reg[142][1]  ( .D(n2382), .CP(clk), .Q(\mem[142][1] ) );
  DFQD1 \mem_reg[142][0]  ( .D(n2381), .CP(clk), .Q(\mem[142][0] ) );
  DFQD1 \mem_reg[143][15]  ( .D(n2380), .CP(clk), .Q(\mem[143][15] ) );
  DFQD1 \mem_reg[143][14]  ( .D(n2379), .CP(clk), .Q(\mem[143][14] ) );
  DFQD1 \mem_reg[143][13]  ( .D(n2378), .CP(clk), .Q(\mem[143][13] ) );
  DFQD1 \mem_reg[143][12]  ( .D(n2377), .CP(clk), .Q(\mem[143][12] ) );
  DFQD1 \mem_reg[143][11]  ( .D(n2376), .CP(clk), .Q(\mem[143][11] ) );
  DFQD1 \mem_reg[143][10]  ( .D(n2375), .CP(clk), .Q(\mem[143][10] ) );
  DFQD1 \mem_reg[143][9]  ( .D(n2374), .CP(clk), .Q(\mem[143][9] ) );
  DFQD1 \mem_reg[143][8]  ( .D(n2373), .CP(clk), .Q(\mem[143][8] ) );
  DFQD1 \mem_reg[143][7]  ( .D(n2372), .CP(clk), .Q(\mem[143][7] ) );
  DFQD1 \mem_reg[143][6]  ( .D(n2371), .CP(clk), .Q(\mem[143][6] ) );
  DFQD1 \mem_reg[143][5]  ( .D(n2370), .CP(clk), .Q(\mem[143][5] ) );
  DFQD1 \mem_reg[143][4]  ( .D(n2369), .CP(clk), .Q(\mem[143][4] ) );
  DFQD1 \mem_reg[143][3]  ( .D(n2368), .CP(clk), .Q(\mem[143][3] ) );
  DFQD1 \mem_reg[143][2]  ( .D(n2367), .CP(clk), .Q(\mem[143][2] ) );
  DFQD1 \mem_reg[143][1]  ( .D(n2366), .CP(clk), .Q(\mem[143][1] ) );
  DFQD1 \mem_reg[143][0]  ( .D(n2365), .CP(clk), .Q(\mem[143][0] ) );
  DFQD1 \mem_reg[144][15]  ( .D(n2364), .CP(clk), .Q(\mem[144][15] ) );
  DFQD1 \mem_reg[144][14]  ( .D(n2363), .CP(clk), .Q(\mem[144][14] ) );
  DFQD1 \mem_reg[144][13]  ( .D(n2362), .CP(clk), .Q(\mem[144][13] ) );
  DFQD1 \mem_reg[144][12]  ( .D(n2361), .CP(clk), .Q(\mem[144][12] ) );
  DFQD1 \mem_reg[144][11]  ( .D(n2360), .CP(clk), .Q(\mem[144][11] ) );
  DFQD1 \mem_reg[144][10]  ( .D(n2359), .CP(clk), .Q(\mem[144][10] ) );
  DFQD1 \mem_reg[144][9]  ( .D(n2358), .CP(clk), .Q(\mem[144][9] ) );
  DFQD1 \mem_reg[144][8]  ( .D(n2357), .CP(clk), .Q(\mem[144][8] ) );
  DFQD1 \mem_reg[144][7]  ( .D(n2356), .CP(clk), .Q(\mem[144][7] ) );
  DFQD1 \mem_reg[144][6]  ( .D(n2355), .CP(clk), .Q(\mem[144][6] ) );
  DFQD1 \mem_reg[144][5]  ( .D(n2354), .CP(clk), .Q(\mem[144][5] ) );
  DFQD1 \mem_reg[144][4]  ( .D(n2353), .CP(clk), .Q(\mem[144][4] ) );
  DFQD1 \mem_reg[144][3]  ( .D(n2352), .CP(clk), .Q(\mem[144][3] ) );
  DFQD1 \mem_reg[144][2]  ( .D(n2351), .CP(clk), .Q(\mem[144][2] ) );
  DFQD1 \mem_reg[144][1]  ( .D(n2350), .CP(clk), .Q(\mem[144][1] ) );
  DFQD1 \mem_reg[144][0]  ( .D(n2349), .CP(clk), .Q(\mem[144][0] ) );
  DFQD1 \mem_reg[145][15]  ( .D(n2348), .CP(clk), .Q(\mem[145][15] ) );
  DFQD1 \mem_reg[145][14]  ( .D(n2347), .CP(clk), .Q(\mem[145][14] ) );
  DFQD1 \mem_reg[145][13]  ( .D(n2346), .CP(clk), .Q(\mem[145][13] ) );
  DFQD1 \mem_reg[145][12]  ( .D(n2345), .CP(clk), .Q(\mem[145][12] ) );
  DFQD1 \mem_reg[145][11]  ( .D(n2344), .CP(clk), .Q(\mem[145][11] ) );
  DFQD1 \mem_reg[145][10]  ( .D(n2343), .CP(clk), .Q(\mem[145][10] ) );
  DFQD1 \mem_reg[145][9]  ( .D(n2342), .CP(clk), .Q(\mem[145][9] ) );
  DFQD1 \mem_reg[145][8]  ( .D(n2341), .CP(clk), .Q(\mem[145][8] ) );
  DFQD1 \mem_reg[145][7]  ( .D(n2340), .CP(clk), .Q(\mem[145][7] ) );
  DFQD1 \mem_reg[145][6]  ( .D(n2339), .CP(clk), .Q(\mem[145][6] ) );
  DFQD1 \mem_reg[145][5]  ( .D(n2338), .CP(clk), .Q(\mem[145][5] ) );
  DFQD1 \mem_reg[145][4]  ( .D(n2337), .CP(clk), .Q(\mem[145][4] ) );
  DFQD1 \mem_reg[145][3]  ( .D(n2336), .CP(clk), .Q(\mem[145][3] ) );
  DFQD1 \mem_reg[145][2]  ( .D(n2335), .CP(clk), .Q(\mem[145][2] ) );
  DFQD1 \mem_reg[145][1]  ( .D(n2334), .CP(clk), .Q(\mem[145][1] ) );
  DFQD1 \mem_reg[145][0]  ( .D(n2333), .CP(clk), .Q(\mem[145][0] ) );
  DFQD1 \mem_reg[146][15]  ( .D(n2332), .CP(clk), .Q(\mem[146][15] ) );
  DFQD1 \mem_reg[146][14]  ( .D(n2331), .CP(clk), .Q(\mem[146][14] ) );
  DFQD1 \mem_reg[146][13]  ( .D(n2330), .CP(clk), .Q(\mem[146][13] ) );
  DFQD1 \mem_reg[146][12]  ( .D(n2329), .CP(clk), .Q(\mem[146][12] ) );
  DFQD1 \mem_reg[146][11]  ( .D(n2328), .CP(clk), .Q(\mem[146][11] ) );
  DFQD1 \mem_reg[146][10]  ( .D(n2327), .CP(clk), .Q(\mem[146][10] ) );
  DFQD1 \mem_reg[146][9]  ( .D(n2326), .CP(clk), .Q(\mem[146][9] ) );
  DFQD1 \mem_reg[146][8]  ( .D(n2325), .CP(clk), .Q(\mem[146][8] ) );
  DFQD1 \mem_reg[146][7]  ( .D(n2324), .CP(clk), .Q(\mem[146][7] ) );
  DFQD1 \mem_reg[146][6]  ( .D(n2323), .CP(clk), .Q(\mem[146][6] ) );
  DFQD1 \mem_reg[146][5]  ( .D(n2322), .CP(clk), .Q(\mem[146][5] ) );
  DFQD1 \mem_reg[146][4]  ( .D(n2321), .CP(clk), .Q(\mem[146][4] ) );
  DFQD1 \mem_reg[146][3]  ( .D(n2320), .CP(clk), .Q(\mem[146][3] ) );
  DFQD1 \mem_reg[146][2]  ( .D(n2319), .CP(clk), .Q(\mem[146][2] ) );
  DFQD1 \mem_reg[146][1]  ( .D(n2318), .CP(clk), .Q(\mem[146][1] ) );
  DFQD1 \mem_reg[146][0]  ( .D(n2317), .CP(clk), .Q(\mem[146][0] ) );
  DFQD1 \mem_reg[147][15]  ( .D(n2316), .CP(clk), .Q(\mem[147][15] ) );
  DFQD1 \mem_reg[147][14]  ( .D(n2315), .CP(clk), .Q(\mem[147][14] ) );
  DFQD1 \mem_reg[147][13]  ( .D(n2314), .CP(clk), .Q(\mem[147][13] ) );
  DFQD1 \mem_reg[147][12]  ( .D(n2313), .CP(clk), .Q(\mem[147][12] ) );
  DFQD1 \mem_reg[147][11]  ( .D(n2312), .CP(clk), .Q(\mem[147][11] ) );
  DFQD1 \mem_reg[147][10]  ( .D(n2311), .CP(clk), .Q(\mem[147][10] ) );
  DFQD1 \mem_reg[147][9]  ( .D(n2310), .CP(clk), .Q(\mem[147][9] ) );
  DFQD1 \mem_reg[147][8]  ( .D(n2309), .CP(clk), .Q(\mem[147][8] ) );
  DFQD1 \mem_reg[147][7]  ( .D(n2308), .CP(clk), .Q(\mem[147][7] ) );
  DFQD1 \mem_reg[147][6]  ( .D(n2307), .CP(clk), .Q(\mem[147][6] ) );
  DFQD1 \mem_reg[147][5]  ( .D(n2306), .CP(clk), .Q(\mem[147][5] ) );
  DFQD1 \mem_reg[147][4]  ( .D(n2305), .CP(clk), .Q(\mem[147][4] ) );
  DFQD1 \mem_reg[147][3]  ( .D(n2304), .CP(clk), .Q(\mem[147][3] ) );
  DFQD1 \mem_reg[147][2]  ( .D(n2303), .CP(clk), .Q(\mem[147][2] ) );
  DFQD1 \mem_reg[147][1]  ( .D(n2302), .CP(clk), .Q(\mem[147][1] ) );
  DFQD1 \mem_reg[147][0]  ( .D(n2301), .CP(clk), .Q(\mem[147][0] ) );
  DFQD1 \mem_reg[148][15]  ( .D(n2300), .CP(clk), .Q(\mem[148][15] ) );
  DFQD1 \mem_reg[148][14]  ( .D(n2299), .CP(clk), .Q(\mem[148][14] ) );
  DFQD1 \mem_reg[148][13]  ( .D(n2298), .CP(clk), .Q(\mem[148][13] ) );
  DFQD1 \mem_reg[148][12]  ( .D(n2297), .CP(clk), .Q(\mem[148][12] ) );
  DFQD1 \mem_reg[148][11]  ( .D(n2296), .CP(clk), .Q(\mem[148][11] ) );
  DFQD1 \mem_reg[148][10]  ( .D(n2295), .CP(clk), .Q(\mem[148][10] ) );
  DFQD1 \mem_reg[148][9]  ( .D(n2294), .CP(clk), .Q(\mem[148][9] ) );
  DFQD1 \mem_reg[148][8]  ( .D(n2293), .CP(clk), .Q(\mem[148][8] ) );
  DFQD1 \mem_reg[148][7]  ( .D(n2292), .CP(clk), .Q(\mem[148][7] ) );
  DFQD1 \mem_reg[148][6]  ( .D(n2291), .CP(clk), .Q(\mem[148][6] ) );
  DFQD1 \mem_reg[148][5]  ( .D(n2290), .CP(clk), .Q(\mem[148][5] ) );
  DFQD1 \mem_reg[148][4]  ( .D(n2289), .CP(clk), .Q(\mem[148][4] ) );
  DFQD1 \mem_reg[148][3]  ( .D(n2288), .CP(clk), .Q(\mem[148][3] ) );
  DFQD1 \mem_reg[148][2]  ( .D(n2287), .CP(clk), .Q(\mem[148][2] ) );
  DFQD1 \mem_reg[148][1]  ( .D(n2286), .CP(clk), .Q(\mem[148][1] ) );
  DFQD1 \mem_reg[148][0]  ( .D(n2285), .CP(clk), .Q(\mem[148][0] ) );
  DFQD1 \mem_reg[149][15]  ( .D(n2284), .CP(clk), .Q(\mem[149][15] ) );
  DFQD1 \mem_reg[149][14]  ( .D(n2283), .CP(clk), .Q(\mem[149][14] ) );
  DFQD1 \mem_reg[149][13]  ( .D(n2282), .CP(clk), .Q(\mem[149][13] ) );
  DFQD1 \mem_reg[149][12]  ( .D(n2281), .CP(clk), .Q(\mem[149][12] ) );
  DFQD1 \mem_reg[149][11]  ( .D(n2280), .CP(clk), .Q(\mem[149][11] ) );
  DFQD1 \mem_reg[149][10]  ( .D(n2279), .CP(clk), .Q(\mem[149][10] ) );
  DFQD1 \mem_reg[149][9]  ( .D(n2278), .CP(clk), .Q(\mem[149][9] ) );
  DFQD1 \mem_reg[149][8]  ( .D(n2277), .CP(clk), .Q(\mem[149][8] ) );
  DFQD1 \mem_reg[149][7]  ( .D(n2276), .CP(clk), .Q(\mem[149][7] ) );
  DFQD1 \mem_reg[149][6]  ( .D(n2275), .CP(clk), .Q(\mem[149][6] ) );
  DFQD1 \mem_reg[149][5]  ( .D(n2274), .CP(clk), .Q(\mem[149][5] ) );
  DFQD1 \mem_reg[149][4]  ( .D(n2273), .CP(clk), .Q(\mem[149][4] ) );
  DFQD1 \mem_reg[149][3]  ( .D(n2272), .CP(clk), .Q(\mem[149][3] ) );
  DFQD1 \mem_reg[149][2]  ( .D(n2271), .CP(clk), .Q(\mem[149][2] ) );
  DFQD1 \mem_reg[149][1]  ( .D(n2270), .CP(clk), .Q(\mem[149][1] ) );
  DFQD1 \mem_reg[149][0]  ( .D(n2269), .CP(clk), .Q(\mem[149][0] ) );
  DFQD1 \mem_reg[150][15]  ( .D(n2268), .CP(clk), .Q(\mem[150][15] ) );
  DFQD1 \mem_reg[150][14]  ( .D(n2267), .CP(clk), .Q(\mem[150][14] ) );
  DFQD1 \mem_reg[150][13]  ( .D(n2266), .CP(clk), .Q(\mem[150][13] ) );
  DFQD1 \mem_reg[150][12]  ( .D(n2265), .CP(clk), .Q(\mem[150][12] ) );
  DFQD1 \mem_reg[150][11]  ( .D(n2264), .CP(clk), .Q(\mem[150][11] ) );
  DFQD1 \mem_reg[150][10]  ( .D(n2263), .CP(clk), .Q(\mem[150][10] ) );
  DFQD1 \mem_reg[150][9]  ( .D(n2262), .CP(clk), .Q(\mem[150][9] ) );
  DFQD1 \mem_reg[150][8]  ( .D(n2261), .CP(clk), .Q(\mem[150][8] ) );
  DFQD1 \mem_reg[150][7]  ( .D(n2260), .CP(clk), .Q(\mem[150][7] ) );
  DFQD1 \mem_reg[150][6]  ( .D(n2259), .CP(clk), .Q(\mem[150][6] ) );
  DFQD1 \mem_reg[150][5]  ( .D(n2258), .CP(clk), .Q(\mem[150][5] ) );
  DFQD1 \mem_reg[150][4]  ( .D(n2257), .CP(clk), .Q(\mem[150][4] ) );
  DFQD1 \mem_reg[150][3]  ( .D(n2256), .CP(clk), .Q(\mem[150][3] ) );
  DFQD1 \mem_reg[150][2]  ( .D(n2255), .CP(clk), .Q(\mem[150][2] ) );
  DFQD1 \mem_reg[150][1]  ( .D(n2254), .CP(clk), .Q(\mem[150][1] ) );
  DFQD1 \mem_reg[150][0]  ( .D(n2253), .CP(clk), .Q(\mem[150][0] ) );
  DFQD1 \mem_reg[151][15]  ( .D(n2252), .CP(clk), .Q(\mem[151][15] ) );
  DFQD1 \mem_reg[151][14]  ( .D(n2251), .CP(clk), .Q(\mem[151][14] ) );
  DFQD1 \mem_reg[151][13]  ( .D(n2250), .CP(clk), .Q(\mem[151][13] ) );
  DFQD1 \mem_reg[151][12]  ( .D(n2249), .CP(clk), .Q(\mem[151][12] ) );
  DFQD1 \mem_reg[151][11]  ( .D(n2248), .CP(clk), .Q(\mem[151][11] ) );
  DFQD1 \mem_reg[151][10]  ( .D(n2247), .CP(clk), .Q(\mem[151][10] ) );
  DFQD1 \mem_reg[151][9]  ( .D(n2246), .CP(clk), .Q(\mem[151][9] ) );
  DFQD1 \mem_reg[151][8]  ( .D(n2245), .CP(clk), .Q(\mem[151][8] ) );
  DFQD1 \mem_reg[151][7]  ( .D(n2244), .CP(clk), .Q(\mem[151][7] ) );
  DFQD1 \mem_reg[151][6]  ( .D(n2243), .CP(clk), .Q(\mem[151][6] ) );
  DFQD1 \mem_reg[151][5]  ( .D(n2242), .CP(clk), .Q(\mem[151][5] ) );
  DFQD1 \mem_reg[151][4]  ( .D(n2241), .CP(clk), .Q(\mem[151][4] ) );
  DFQD1 \mem_reg[151][3]  ( .D(n2240), .CP(clk), .Q(\mem[151][3] ) );
  DFQD1 \mem_reg[151][2]  ( .D(n2239), .CP(clk), .Q(\mem[151][2] ) );
  DFQD1 \mem_reg[151][1]  ( .D(n2238), .CP(clk), .Q(\mem[151][1] ) );
  DFQD1 \mem_reg[151][0]  ( .D(n2237), .CP(clk), .Q(\mem[151][0] ) );
  DFQD1 \mem_reg[152][15]  ( .D(n2236), .CP(clk), .Q(\mem[152][15] ) );
  DFQD1 \mem_reg[152][14]  ( .D(n2235), .CP(clk), .Q(\mem[152][14] ) );
  DFQD1 \mem_reg[152][13]  ( .D(n2234), .CP(clk), .Q(\mem[152][13] ) );
  DFQD1 \mem_reg[152][12]  ( .D(n2233), .CP(clk), .Q(\mem[152][12] ) );
  DFQD1 \mem_reg[152][11]  ( .D(n2232), .CP(clk), .Q(\mem[152][11] ) );
  DFQD1 \mem_reg[152][10]  ( .D(n2231), .CP(clk), .Q(\mem[152][10] ) );
  DFQD1 \mem_reg[152][9]  ( .D(n2230), .CP(clk), .Q(\mem[152][9] ) );
  DFQD1 \mem_reg[152][8]  ( .D(n2229), .CP(clk), .Q(\mem[152][8] ) );
  DFQD1 \mem_reg[152][7]  ( .D(n2228), .CP(clk), .Q(\mem[152][7] ) );
  DFQD1 \mem_reg[152][6]  ( .D(n2227), .CP(clk), .Q(\mem[152][6] ) );
  DFQD1 \mem_reg[152][5]  ( .D(n2226), .CP(clk), .Q(\mem[152][5] ) );
  DFQD1 \mem_reg[152][4]  ( .D(n2225), .CP(clk), .Q(\mem[152][4] ) );
  DFQD1 \mem_reg[152][3]  ( .D(n2224), .CP(clk), .Q(\mem[152][3] ) );
  DFQD1 \mem_reg[152][2]  ( .D(n2223), .CP(clk), .Q(\mem[152][2] ) );
  DFQD1 \mem_reg[152][1]  ( .D(n2222), .CP(clk), .Q(\mem[152][1] ) );
  DFQD1 \mem_reg[152][0]  ( .D(n2221), .CP(clk), .Q(\mem[152][0] ) );
  DFQD1 \mem_reg[153][15]  ( .D(n2220), .CP(clk), .Q(\mem[153][15] ) );
  DFQD1 \mem_reg[153][14]  ( .D(n2219), .CP(clk), .Q(\mem[153][14] ) );
  DFQD1 \mem_reg[153][13]  ( .D(n2218), .CP(clk), .Q(\mem[153][13] ) );
  DFQD1 \mem_reg[153][12]  ( .D(n2217), .CP(clk), .Q(\mem[153][12] ) );
  DFQD1 \mem_reg[153][11]  ( .D(n2216), .CP(clk), .Q(\mem[153][11] ) );
  DFQD1 \mem_reg[153][10]  ( .D(n2215), .CP(clk), .Q(\mem[153][10] ) );
  DFQD1 \mem_reg[153][9]  ( .D(n2214), .CP(clk), .Q(\mem[153][9] ) );
  DFQD1 \mem_reg[153][8]  ( .D(n2213), .CP(clk), .Q(\mem[153][8] ) );
  DFQD1 \mem_reg[153][7]  ( .D(n2212), .CP(clk), .Q(\mem[153][7] ) );
  DFQD1 \mem_reg[153][6]  ( .D(n2211), .CP(clk), .Q(\mem[153][6] ) );
  DFQD1 \mem_reg[153][5]  ( .D(n2210), .CP(clk), .Q(\mem[153][5] ) );
  DFQD1 \mem_reg[153][4]  ( .D(n2209), .CP(clk), .Q(\mem[153][4] ) );
  DFQD1 \mem_reg[153][3]  ( .D(n2208), .CP(clk), .Q(\mem[153][3] ) );
  DFQD1 \mem_reg[153][2]  ( .D(n2207), .CP(clk), .Q(\mem[153][2] ) );
  DFQD1 \mem_reg[153][1]  ( .D(n2206), .CP(clk), .Q(\mem[153][1] ) );
  DFQD1 \mem_reg[153][0]  ( .D(n2205), .CP(clk), .Q(\mem[153][0] ) );
  DFQD1 \mem_reg[154][15]  ( .D(n2204), .CP(clk), .Q(\mem[154][15] ) );
  DFQD1 \mem_reg[154][14]  ( .D(n2203), .CP(clk), .Q(\mem[154][14] ) );
  DFQD1 \mem_reg[154][13]  ( .D(n2202), .CP(clk), .Q(\mem[154][13] ) );
  DFQD1 \mem_reg[154][12]  ( .D(n2201), .CP(clk), .Q(\mem[154][12] ) );
  DFQD1 \mem_reg[154][11]  ( .D(n2200), .CP(clk), .Q(\mem[154][11] ) );
  DFQD1 \mem_reg[154][10]  ( .D(n2199), .CP(clk), .Q(\mem[154][10] ) );
  DFQD1 \mem_reg[154][9]  ( .D(n2198), .CP(clk), .Q(\mem[154][9] ) );
  DFQD1 \mem_reg[154][8]  ( .D(n2197), .CP(clk), .Q(\mem[154][8] ) );
  DFQD1 \mem_reg[154][7]  ( .D(n2196), .CP(clk), .Q(\mem[154][7] ) );
  DFQD1 \mem_reg[154][6]  ( .D(n2195), .CP(clk), .Q(\mem[154][6] ) );
  DFQD1 \mem_reg[154][5]  ( .D(n2194), .CP(clk), .Q(\mem[154][5] ) );
  DFQD1 \mem_reg[154][4]  ( .D(n2193), .CP(clk), .Q(\mem[154][4] ) );
  DFQD1 \mem_reg[154][3]  ( .D(n2192), .CP(clk), .Q(\mem[154][3] ) );
  DFQD1 \mem_reg[154][2]  ( .D(n2191), .CP(clk), .Q(\mem[154][2] ) );
  DFQD1 \mem_reg[154][1]  ( .D(n2190), .CP(clk), .Q(\mem[154][1] ) );
  DFQD1 \mem_reg[154][0]  ( .D(n2189), .CP(clk), .Q(\mem[154][0] ) );
  DFQD1 \mem_reg[155][15]  ( .D(n2188), .CP(clk), .Q(\mem[155][15] ) );
  DFQD1 \mem_reg[155][14]  ( .D(n2187), .CP(clk), .Q(\mem[155][14] ) );
  DFQD1 \mem_reg[155][13]  ( .D(n2186), .CP(clk), .Q(\mem[155][13] ) );
  DFQD1 \mem_reg[155][12]  ( .D(n2185), .CP(clk), .Q(\mem[155][12] ) );
  DFQD1 \mem_reg[155][11]  ( .D(n2184), .CP(clk), .Q(\mem[155][11] ) );
  DFQD1 \mem_reg[155][10]  ( .D(n2183), .CP(clk), .Q(\mem[155][10] ) );
  DFQD1 \mem_reg[155][9]  ( .D(n2182), .CP(clk), .Q(\mem[155][9] ) );
  DFQD1 \mem_reg[155][8]  ( .D(n2181), .CP(clk), .Q(\mem[155][8] ) );
  DFQD1 \mem_reg[155][7]  ( .D(n2180), .CP(clk), .Q(\mem[155][7] ) );
  DFQD1 \mem_reg[155][6]  ( .D(n2179), .CP(clk), .Q(\mem[155][6] ) );
  DFQD1 \mem_reg[155][5]  ( .D(n2178), .CP(clk), .Q(\mem[155][5] ) );
  DFQD1 \mem_reg[155][4]  ( .D(n2177), .CP(clk), .Q(\mem[155][4] ) );
  DFQD1 \mem_reg[155][3]  ( .D(n2176), .CP(clk), .Q(\mem[155][3] ) );
  DFQD1 \mem_reg[155][2]  ( .D(n2175), .CP(clk), .Q(\mem[155][2] ) );
  DFQD1 \mem_reg[155][1]  ( .D(n2174), .CP(clk), .Q(\mem[155][1] ) );
  DFQD1 \mem_reg[155][0]  ( .D(n2173), .CP(clk), .Q(\mem[155][0] ) );
  DFQD1 \mem_reg[156][15]  ( .D(n2172), .CP(clk), .Q(\mem[156][15] ) );
  DFQD1 \mem_reg[156][14]  ( .D(n2171), .CP(clk), .Q(\mem[156][14] ) );
  DFQD1 \mem_reg[156][13]  ( .D(n2170), .CP(clk), .Q(\mem[156][13] ) );
  DFQD1 \mem_reg[156][12]  ( .D(n2169), .CP(clk), .Q(\mem[156][12] ) );
  DFQD1 \mem_reg[156][11]  ( .D(n2168), .CP(clk), .Q(\mem[156][11] ) );
  DFQD1 \mem_reg[156][10]  ( .D(n2167), .CP(clk), .Q(\mem[156][10] ) );
  DFQD1 \mem_reg[156][9]  ( .D(n2166), .CP(clk), .Q(\mem[156][9] ) );
  DFQD1 \mem_reg[156][8]  ( .D(n2165), .CP(clk), .Q(\mem[156][8] ) );
  DFQD1 \mem_reg[156][7]  ( .D(n2164), .CP(clk), .Q(\mem[156][7] ) );
  DFQD1 \mem_reg[156][6]  ( .D(n2163), .CP(clk), .Q(\mem[156][6] ) );
  DFQD1 \mem_reg[156][5]  ( .D(n2162), .CP(clk), .Q(\mem[156][5] ) );
  DFQD1 \mem_reg[156][4]  ( .D(n2161), .CP(clk), .Q(\mem[156][4] ) );
  DFQD1 \mem_reg[156][3]  ( .D(n2160), .CP(clk), .Q(\mem[156][3] ) );
  DFQD1 \mem_reg[156][2]  ( .D(n2159), .CP(clk), .Q(\mem[156][2] ) );
  DFQD1 \mem_reg[156][1]  ( .D(n2158), .CP(clk), .Q(\mem[156][1] ) );
  DFQD1 \mem_reg[156][0]  ( .D(n2157), .CP(clk), .Q(\mem[156][0] ) );
  DFQD1 \mem_reg[157][15]  ( .D(n2156), .CP(clk), .Q(\mem[157][15] ) );
  DFQD1 \mem_reg[157][14]  ( .D(n2155), .CP(clk), .Q(\mem[157][14] ) );
  DFQD1 \mem_reg[157][13]  ( .D(n2154), .CP(clk), .Q(\mem[157][13] ) );
  DFQD1 \mem_reg[157][12]  ( .D(n2153), .CP(clk), .Q(\mem[157][12] ) );
  DFQD1 \mem_reg[157][11]  ( .D(n2152), .CP(clk), .Q(\mem[157][11] ) );
  DFQD1 \mem_reg[157][10]  ( .D(n2151), .CP(clk), .Q(\mem[157][10] ) );
  DFQD1 \mem_reg[157][9]  ( .D(n2150), .CP(clk), .Q(\mem[157][9] ) );
  DFQD1 \mem_reg[157][8]  ( .D(n2149), .CP(clk), .Q(\mem[157][8] ) );
  DFQD1 \mem_reg[157][7]  ( .D(n2148), .CP(clk), .Q(\mem[157][7] ) );
  DFQD1 \mem_reg[157][6]  ( .D(n2147), .CP(clk), .Q(\mem[157][6] ) );
  DFQD1 \mem_reg[157][5]  ( .D(n2146), .CP(clk), .Q(\mem[157][5] ) );
  DFQD1 \mem_reg[157][4]  ( .D(n2145), .CP(clk), .Q(\mem[157][4] ) );
  DFQD1 \mem_reg[157][3]  ( .D(n2144), .CP(clk), .Q(\mem[157][3] ) );
  DFQD1 \mem_reg[157][2]  ( .D(n2143), .CP(clk), .Q(\mem[157][2] ) );
  DFQD1 \mem_reg[157][1]  ( .D(n2142), .CP(clk), .Q(\mem[157][1] ) );
  DFQD1 \mem_reg[157][0]  ( .D(n2141), .CP(clk), .Q(\mem[157][0] ) );
  DFQD1 \mem_reg[158][15]  ( .D(n2140), .CP(clk), .Q(\mem[158][15] ) );
  DFQD1 \mem_reg[158][14]  ( .D(n2139), .CP(clk), .Q(\mem[158][14] ) );
  DFQD1 \mem_reg[158][13]  ( .D(n2138), .CP(clk), .Q(\mem[158][13] ) );
  DFQD1 \mem_reg[158][12]  ( .D(n2137), .CP(clk), .Q(\mem[158][12] ) );
  DFQD1 \mem_reg[158][11]  ( .D(n2136), .CP(clk), .Q(\mem[158][11] ) );
  DFQD1 \mem_reg[158][10]  ( .D(n2135), .CP(clk), .Q(\mem[158][10] ) );
  DFQD1 \mem_reg[158][9]  ( .D(n2134), .CP(clk), .Q(\mem[158][9] ) );
  DFQD1 \mem_reg[158][8]  ( .D(n2133), .CP(clk), .Q(\mem[158][8] ) );
  DFQD1 \mem_reg[158][7]  ( .D(n2132), .CP(clk), .Q(\mem[158][7] ) );
  DFQD1 \mem_reg[158][6]  ( .D(n2131), .CP(clk), .Q(\mem[158][6] ) );
  DFQD1 \mem_reg[158][5]  ( .D(n2130), .CP(clk), .Q(\mem[158][5] ) );
  DFQD1 \mem_reg[158][4]  ( .D(n2129), .CP(clk), .Q(\mem[158][4] ) );
  DFQD1 \mem_reg[158][3]  ( .D(n2128), .CP(clk), .Q(\mem[158][3] ) );
  DFQD1 \mem_reg[158][2]  ( .D(n2127), .CP(clk), .Q(\mem[158][2] ) );
  DFQD1 \mem_reg[158][1]  ( .D(n2126), .CP(clk), .Q(\mem[158][1] ) );
  DFQD1 \mem_reg[158][0]  ( .D(n2125), .CP(clk), .Q(\mem[158][0] ) );
  DFQD1 \mem_reg[159][15]  ( .D(n2124), .CP(clk), .Q(\mem[159][15] ) );
  DFQD1 \mem_reg[159][14]  ( .D(n2123), .CP(clk), .Q(\mem[159][14] ) );
  DFQD1 \mem_reg[159][13]  ( .D(n2122), .CP(clk), .Q(\mem[159][13] ) );
  DFQD1 \mem_reg[159][12]  ( .D(n2121), .CP(clk), .Q(\mem[159][12] ) );
  DFQD1 \mem_reg[159][11]  ( .D(n2120), .CP(clk), .Q(\mem[159][11] ) );
  DFQD1 \mem_reg[159][10]  ( .D(n2119), .CP(clk), .Q(\mem[159][10] ) );
  DFQD1 \mem_reg[159][9]  ( .D(n2118), .CP(clk), .Q(\mem[159][9] ) );
  DFQD1 \mem_reg[159][8]  ( .D(n2117), .CP(clk), .Q(\mem[159][8] ) );
  DFQD1 \mem_reg[159][7]  ( .D(n2116), .CP(clk), .Q(\mem[159][7] ) );
  DFQD1 \mem_reg[159][6]  ( .D(n2115), .CP(clk), .Q(\mem[159][6] ) );
  DFQD1 \mem_reg[159][5]  ( .D(n2114), .CP(clk), .Q(\mem[159][5] ) );
  DFQD1 \mem_reg[159][4]  ( .D(n2113), .CP(clk), .Q(\mem[159][4] ) );
  DFQD1 \mem_reg[159][3]  ( .D(n2112), .CP(clk), .Q(\mem[159][3] ) );
  DFQD1 \mem_reg[159][2]  ( .D(n2111), .CP(clk), .Q(\mem[159][2] ) );
  DFQD1 \mem_reg[159][1]  ( .D(n2110), .CP(clk), .Q(\mem[159][1] ) );
  DFQD1 \mem_reg[159][0]  ( .D(n2109), .CP(clk), .Q(\mem[159][0] ) );
  DFQD1 \mem_reg[160][15]  ( .D(n2108), .CP(clk), .Q(\mem[160][15] ) );
  DFQD1 \mem_reg[160][14]  ( .D(n2107), .CP(clk), .Q(\mem[160][14] ) );
  DFQD1 \mem_reg[160][13]  ( .D(n2106), .CP(clk), .Q(\mem[160][13] ) );
  DFQD1 \mem_reg[160][12]  ( .D(n2105), .CP(clk), .Q(\mem[160][12] ) );
  DFQD1 \mem_reg[160][11]  ( .D(n2104), .CP(clk), .Q(\mem[160][11] ) );
  DFQD1 \mem_reg[160][10]  ( .D(n2103), .CP(clk), .Q(\mem[160][10] ) );
  DFQD1 \mem_reg[160][9]  ( .D(n2102), .CP(clk), .Q(\mem[160][9] ) );
  DFQD1 \mem_reg[160][8]  ( .D(n2101), .CP(clk), .Q(\mem[160][8] ) );
  DFQD1 \mem_reg[160][7]  ( .D(n2100), .CP(clk), .Q(\mem[160][7] ) );
  DFQD1 \mem_reg[160][6]  ( .D(n2099), .CP(clk), .Q(\mem[160][6] ) );
  DFQD1 \mem_reg[160][5]  ( .D(n2098), .CP(clk), .Q(\mem[160][5] ) );
  DFQD1 \mem_reg[160][4]  ( .D(n2097), .CP(clk), .Q(\mem[160][4] ) );
  DFQD1 \mem_reg[160][3]  ( .D(n2096), .CP(clk), .Q(\mem[160][3] ) );
  DFQD1 \mem_reg[160][2]  ( .D(n2095), .CP(clk), .Q(\mem[160][2] ) );
  DFQD1 \mem_reg[160][1]  ( .D(n2094), .CP(clk), .Q(\mem[160][1] ) );
  DFQD1 \mem_reg[160][0]  ( .D(n2093), .CP(clk), .Q(\mem[160][0] ) );
  DFQD1 \mem_reg[161][15]  ( .D(n2092), .CP(clk), .Q(\mem[161][15] ) );
  DFQD1 \mem_reg[161][14]  ( .D(n2091), .CP(clk), .Q(\mem[161][14] ) );
  DFQD1 \mem_reg[161][13]  ( .D(n2090), .CP(clk), .Q(\mem[161][13] ) );
  DFQD1 \mem_reg[161][12]  ( .D(n2089), .CP(clk), .Q(\mem[161][12] ) );
  DFQD1 \mem_reg[161][11]  ( .D(n2088), .CP(clk), .Q(\mem[161][11] ) );
  DFQD1 \mem_reg[161][10]  ( .D(n2087), .CP(clk), .Q(\mem[161][10] ) );
  DFQD1 \mem_reg[161][9]  ( .D(n2086), .CP(clk), .Q(\mem[161][9] ) );
  DFQD1 \mem_reg[161][8]  ( .D(n2085), .CP(clk), .Q(\mem[161][8] ) );
  DFQD1 \mem_reg[161][7]  ( .D(n2084), .CP(clk), .Q(\mem[161][7] ) );
  DFQD1 \mem_reg[161][6]  ( .D(n2083), .CP(clk), .Q(\mem[161][6] ) );
  DFQD1 \mem_reg[161][5]  ( .D(n2082), .CP(clk), .Q(\mem[161][5] ) );
  DFQD1 \mem_reg[161][4]  ( .D(n2081), .CP(clk), .Q(\mem[161][4] ) );
  DFQD1 \mem_reg[161][3]  ( .D(n2080), .CP(clk), .Q(\mem[161][3] ) );
  DFQD1 \mem_reg[161][2]  ( .D(n2079), .CP(clk), .Q(\mem[161][2] ) );
  DFQD1 \mem_reg[161][1]  ( .D(n2078), .CP(clk), .Q(\mem[161][1] ) );
  DFQD1 \mem_reg[161][0]  ( .D(n2077), .CP(clk), .Q(\mem[161][0] ) );
  DFQD1 \mem_reg[162][15]  ( .D(n2076), .CP(clk), .Q(\mem[162][15] ) );
  DFQD1 \mem_reg[162][14]  ( .D(n2075), .CP(clk), .Q(\mem[162][14] ) );
  DFQD1 \mem_reg[162][13]  ( .D(n2074), .CP(clk), .Q(\mem[162][13] ) );
  DFQD1 \mem_reg[162][12]  ( .D(n2073), .CP(clk), .Q(\mem[162][12] ) );
  DFQD1 \mem_reg[162][11]  ( .D(n2072), .CP(clk), .Q(\mem[162][11] ) );
  DFQD1 \mem_reg[162][10]  ( .D(n2071), .CP(clk), .Q(\mem[162][10] ) );
  DFQD1 \mem_reg[162][9]  ( .D(n2070), .CP(clk), .Q(\mem[162][9] ) );
  DFQD1 \mem_reg[162][8]  ( .D(n2069), .CP(clk), .Q(\mem[162][8] ) );
  DFQD1 \mem_reg[162][7]  ( .D(n2068), .CP(clk), .Q(\mem[162][7] ) );
  DFQD1 \mem_reg[162][6]  ( .D(n2067), .CP(clk), .Q(\mem[162][6] ) );
  DFQD1 \mem_reg[162][5]  ( .D(n2066), .CP(clk), .Q(\mem[162][5] ) );
  DFQD1 \mem_reg[162][4]  ( .D(n2065), .CP(clk), .Q(\mem[162][4] ) );
  DFQD1 \mem_reg[162][3]  ( .D(n2064), .CP(clk), .Q(\mem[162][3] ) );
  DFQD1 \mem_reg[162][2]  ( .D(n2063), .CP(clk), .Q(\mem[162][2] ) );
  DFQD1 \mem_reg[162][1]  ( .D(n2062), .CP(clk), .Q(\mem[162][1] ) );
  DFQD1 \mem_reg[162][0]  ( .D(n2061), .CP(clk), .Q(\mem[162][0] ) );
  DFQD1 \mem_reg[163][15]  ( .D(n2060), .CP(clk), .Q(\mem[163][15] ) );
  DFQD1 \mem_reg[163][14]  ( .D(n2059), .CP(clk), .Q(\mem[163][14] ) );
  DFQD1 \mem_reg[163][13]  ( .D(n2058), .CP(clk), .Q(\mem[163][13] ) );
  DFQD1 \mem_reg[163][12]  ( .D(n2057), .CP(clk), .Q(\mem[163][12] ) );
  DFQD1 \mem_reg[163][11]  ( .D(n2056), .CP(clk), .Q(\mem[163][11] ) );
  DFQD1 \mem_reg[163][10]  ( .D(n2055), .CP(clk), .Q(\mem[163][10] ) );
  DFQD1 \mem_reg[163][9]  ( .D(n2054), .CP(clk), .Q(\mem[163][9] ) );
  DFQD1 \mem_reg[163][8]  ( .D(n2053), .CP(clk), .Q(\mem[163][8] ) );
  DFQD1 \mem_reg[163][7]  ( .D(n2052), .CP(clk), .Q(\mem[163][7] ) );
  DFQD1 \mem_reg[163][6]  ( .D(n2051), .CP(clk), .Q(\mem[163][6] ) );
  DFQD1 \mem_reg[163][5]  ( .D(n2050), .CP(clk), .Q(\mem[163][5] ) );
  DFQD1 \mem_reg[163][4]  ( .D(n2049), .CP(clk), .Q(\mem[163][4] ) );
  DFQD1 \mem_reg[163][3]  ( .D(n2048), .CP(clk), .Q(\mem[163][3] ) );
  DFQD1 \mem_reg[163][2]  ( .D(n2047), .CP(clk), .Q(\mem[163][2] ) );
  DFQD1 \mem_reg[163][1]  ( .D(n2046), .CP(clk), .Q(\mem[163][1] ) );
  DFQD1 \mem_reg[163][0]  ( .D(n2045), .CP(clk), .Q(\mem[163][0] ) );
  DFQD1 \mem_reg[164][15]  ( .D(n2044), .CP(clk), .Q(\mem[164][15] ) );
  DFQD1 \mem_reg[164][14]  ( .D(n2043), .CP(clk), .Q(\mem[164][14] ) );
  DFQD1 \mem_reg[164][13]  ( .D(n2042), .CP(clk), .Q(\mem[164][13] ) );
  DFQD1 \mem_reg[164][12]  ( .D(n2041), .CP(clk), .Q(\mem[164][12] ) );
  DFQD1 \mem_reg[164][11]  ( .D(n2040), .CP(clk), .Q(\mem[164][11] ) );
  DFQD1 \mem_reg[164][10]  ( .D(n2039), .CP(clk), .Q(\mem[164][10] ) );
  DFQD1 \mem_reg[164][9]  ( .D(n2038), .CP(clk), .Q(\mem[164][9] ) );
  DFQD1 \mem_reg[164][8]  ( .D(n2037), .CP(clk), .Q(\mem[164][8] ) );
  DFQD1 \mem_reg[164][7]  ( .D(n2036), .CP(clk), .Q(\mem[164][7] ) );
  DFQD1 \mem_reg[164][6]  ( .D(n2035), .CP(clk), .Q(\mem[164][6] ) );
  DFQD1 \mem_reg[164][5]  ( .D(n2034), .CP(clk), .Q(\mem[164][5] ) );
  DFQD1 \mem_reg[164][4]  ( .D(n2033), .CP(clk), .Q(\mem[164][4] ) );
  DFQD1 \mem_reg[164][3]  ( .D(n2032), .CP(clk), .Q(\mem[164][3] ) );
  DFQD1 \mem_reg[164][2]  ( .D(n2031), .CP(clk), .Q(\mem[164][2] ) );
  DFQD1 \mem_reg[164][1]  ( .D(n2030), .CP(clk), .Q(\mem[164][1] ) );
  DFQD1 \mem_reg[164][0]  ( .D(n2029), .CP(clk), .Q(\mem[164][0] ) );
  DFQD1 \mem_reg[165][15]  ( .D(n2028), .CP(clk), .Q(\mem[165][15] ) );
  DFQD1 \mem_reg[165][14]  ( .D(n2027), .CP(clk), .Q(\mem[165][14] ) );
  DFQD1 \mem_reg[165][13]  ( .D(n2026), .CP(clk), .Q(\mem[165][13] ) );
  DFQD1 \mem_reg[165][12]  ( .D(n2025), .CP(clk), .Q(\mem[165][12] ) );
  DFQD1 \mem_reg[165][11]  ( .D(n2024), .CP(clk), .Q(\mem[165][11] ) );
  DFQD1 \mem_reg[165][10]  ( .D(n2023), .CP(clk), .Q(\mem[165][10] ) );
  DFQD1 \mem_reg[165][9]  ( .D(n2022), .CP(clk), .Q(\mem[165][9] ) );
  DFQD1 \mem_reg[165][8]  ( .D(n2021), .CP(clk), .Q(\mem[165][8] ) );
  DFQD1 \mem_reg[165][7]  ( .D(n2020), .CP(clk), .Q(\mem[165][7] ) );
  DFQD1 \mem_reg[165][6]  ( .D(n2019), .CP(clk), .Q(\mem[165][6] ) );
  DFQD1 \mem_reg[165][5]  ( .D(n2018), .CP(clk), .Q(\mem[165][5] ) );
  DFQD1 \mem_reg[165][4]  ( .D(n2017), .CP(clk), .Q(\mem[165][4] ) );
  DFQD1 \mem_reg[165][3]  ( .D(n2016), .CP(clk), .Q(\mem[165][3] ) );
  DFQD1 \mem_reg[165][2]  ( .D(n2015), .CP(clk), .Q(\mem[165][2] ) );
  DFQD1 \mem_reg[165][1]  ( .D(n2014), .CP(clk), .Q(\mem[165][1] ) );
  DFQD1 \mem_reg[165][0]  ( .D(n2013), .CP(clk), .Q(\mem[165][0] ) );
  DFQD1 \mem_reg[166][15]  ( .D(n2012), .CP(clk), .Q(\mem[166][15] ) );
  DFQD1 \mem_reg[166][14]  ( .D(n2011), .CP(clk), .Q(\mem[166][14] ) );
  DFQD1 \mem_reg[166][13]  ( .D(n2010), .CP(clk), .Q(\mem[166][13] ) );
  DFQD1 \mem_reg[166][12]  ( .D(n2009), .CP(clk), .Q(\mem[166][12] ) );
  DFQD1 \mem_reg[166][11]  ( .D(n2008), .CP(clk), .Q(\mem[166][11] ) );
  DFQD1 \mem_reg[166][10]  ( .D(n2007), .CP(clk), .Q(\mem[166][10] ) );
  DFQD1 \mem_reg[166][9]  ( .D(n2006), .CP(clk), .Q(\mem[166][9] ) );
  DFQD1 \mem_reg[166][8]  ( .D(n2005), .CP(clk), .Q(\mem[166][8] ) );
  DFQD1 \mem_reg[166][7]  ( .D(n2004), .CP(clk), .Q(\mem[166][7] ) );
  DFQD1 \mem_reg[166][6]  ( .D(n2003), .CP(clk), .Q(\mem[166][6] ) );
  DFQD1 \mem_reg[166][5]  ( .D(n2002), .CP(clk), .Q(\mem[166][5] ) );
  DFQD1 \mem_reg[166][4]  ( .D(n2001), .CP(clk), .Q(\mem[166][4] ) );
  DFQD1 \mem_reg[166][3]  ( .D(n2000), .CP(clk), .Q(\mem[166][3] ) );
  DFQD1 \mem_reg[166][2]  ( .D(n1999), .CP(clk), .Q(\mem[166][2] ) );
  DFQD1 \mem_reg[166][1]  ( .D(n1998), .CP(clk), .Q(\mem[166][1] ) );
  DFQD1 \mem_reg[166][0]  ( .D(n1997), .CP(clk), .Q(\mem[166][0] ) );
  DFQD1 \mem_reg[167][15]  ( .D(n1996), .CP(clk), .Q(\mem[167][15] ) );
  DFQD1 \mem_reg[167][14]  ( .D(n1995), .CP(clk), .Q(\mem[167][14] ) );
  DFQD1 \mem_reg[167][13]  ( .D(n1994), .CP(clk), .Q(\mem[167][13] ) );
  DFQD1 \mem_reg[167][12]  ( .D(n1993), .CP(clk), .Q(\mem[167][12] ) );
  DFQD1 \mem_reg[167][11]  ( .D(n1992), .CP(clk), .Q(\mem[167][11] ) );
  DFQD1 \mem_reg[167][10]  ( .D(n1991), .CP(clk), .Q(\mem[167][10] ) );
  DFQD1 \mem_reg[167][9]  ( .D(n1990), .CP(clk), .Q(\mem[167][9] ) );
  DFQD1 \mem_reg[167][8]  ( .D(n1989), .CP(clk), .Q(\mem[167][8] ) );
  DFQD1 \mem_reg[167][7]  ( .D(n1988), .CP(clk), .Q(\mem[167][7] ) );
  DFQD1 \mem_reg[167][6]  ( .D(n1987), .CP(clk), .Q(\mem[167][6] ) );
  DFQD1 \mem_reg[167][5]  ( .D(n1986), .CP(clk), .Q(\mem[167][5] ) );
  DFQD1 \mem_reg[167][4]  ( .D(n1985), .CP(clk), .Q(\mem[167][4] ) );
  DFQD1 \mem_reg[167][3]  ( .D(n1984), .CP(clk), .Q(\mem[167][3] ) );
  DFQD1 \mem_reg[167][2]  ( .D(n1983), .CP(clk), .Q(\mem[167][2] ) );
  DFQD1 \mem_reg[167][1]  ( .D(n1982), .CP(clk), .Q(\mem[167][1] ) );
  DFQD1 \mem_reg[167][0]  ( .D(n1981), .CP(clk), .Q(\mem[167][0] ) );
  DFQD1 \mem_reg[168][15]  ( .D(n1980), .CP(clk), .Q(\mem[168][15] ) );
  DFQD1 \mem_reg[168][14]  ( .D(n1979), .CP(clk), .Q(\mem[168][14] ) );
  DFQD1 \mem_reg[168][13]  ( .D(n1978), .CP(clk), .Q(\mem[168][13] ) );
  DFQD1 \mem_reg[168][12]  ( .D(n1977), .CP(clk), .Q(\mem[168][12] ) );
  DFQD1 \mem_reg[168][11]  ( .D(n1976), .CP(clk), .Q(\mem[168][11] ) );
  DFQD1 \mem_reg[168][10]  ( .D(n1975), .CP(clk), .Q(\mem[168][10] ) );
  DFQD1 \mem_reg[168][9]  ( .D(n1974), .CP(clk), .Q(\mem[168][9] ) );
  DFQD1 \mem_reg[168][8]  ( .D(n1973), .CP(clk), .Q(\mem[168][8] ) );
  DFQD1 \mem_reg[168][7]  ( .D(n1972), .CP(clk), .Q(\mem[168][7] ) );
  DFQD1 \mem_reg[168][6]  ( .D(n1971), .CP(clk), .Q(\mem[168][6] ) );
  DFQD1 \mem_reg[168][5]  ( .D(n1970), .CP(clk), .Q(\mem[168][5] ) );
  DFQD1 \mem_reg[168][4]  ( .D(n1969), .CP(clk), .Q(\mem[168][4] ) );
  DFQD1 \mem_reg[168][3]  ( .D(n1968), .CP(clk), .Q(\mem[168][3] ) );
  DFQD1 \mem_reg[168][2]  ( .D(n1967), .CP(clk), .Q(\mem[168][2] ) );
  DFQD1 \mem_reg[168][1]  ( .D(n1966), .CP(clk), .Q(\mem[168][1] ) );
  DFQD1 \mem_reg[168][0]  ( .D(n1965), .CP(clk), .Q(\mem[168][0] ) );
  DFQD1 \mem_reg[169][15]  ( .D(n1964), .CP(clk), .Q(\mem[169][15] ) );
  DFQD1 \mem_reg[169][14]  ( .D(n1963), .CP(clk), .Q(\mem[169][14] ) );
  DFQD1 \mem_reg[169][13]  ( .D(n1962), .CP(clk), .Q(\mem[169][13] ) );
  DFQD1 \mem_reg[169][12]  ( .D(n1961), .CP(clk), .Q(\mem[169][12] ) );
  DFQD1 \mem_reg[169][11]  ( .D(n1960), .CP(clk), .Q(\mem[169][11] ) );
  DFQD1 \mem_reg[169][10]  ( .D(n1959), .CP(clk), .Q(\mem[169][10] ) );
  DFQD1 \mem_reg[169][9]  ( .D(n1958), .CP(clk), .Q(\mem[169][9] ) );
  DFQD1 \mem_reg[169][8]  ( .D(n1957), .CP(clk), .Q(\mem[169][8] ) );
  DFQD1 \mem_reg[169][7]  ( .D(n1956), .CP(clk), .Q(\mem[169][7] ) );
  DFQD1 \mem_reg[169][6]  ( .D(n1955), .CP(clk), .Q(\mem[169][6] ) );
  DFQD1 \mem_reg[169][5]  ( .D(n1954), .CP(clk), .Q(\mem[169][5] ) );
  DFQD1 \mem_reg[169][4]  ( .D(n1953), .CP(clk), .Q(\mem[169][4] ) );
  DFQD1 \mem_reg[169][3]  ( .D(n1952), .CP(clk), .Q(\mem[169][3] ) );
  DFQD1 \mem_reg[169][2]  ( .D(n1951), .CP(clk), .Q(\mem[169][2] ) );
  DFQD1 \mem_reg[169][1]  ( .D(n1950), .CP(clk), .Q(\mem[169][1] ) );
  DFQD1 \mem_reg[169][0]  ( .D(n1949), .CP(clk), .Q(\mem[169][0] ) );
  DFQD1 \mem_reg[170][15]  ( .D(n1948), .CP(clk), .Q(\mem[170][15] ) );
  DFQD1 \mem_reg[170][14]  ( .D(n1947), .CP(clk), .Q(\mem[170][14] ) );
  DFQD1 \mem_reg[170][13]  ( .D(n1946), .CP(clk), .Q(\mem[170][13] ) );
  DFQD1 \mem_reg[170][12]  ( .D(n1945), .CP(clk), .Q(\mem[170][12] ) );
  DFQD1 \mem_reg[170][11]  ( .D(n1944), .CP(clk), .Q(\mem[170][11] ) );
  DFQD1 \mem_reg[170][10]  ( .D(n1943), .CP(clk), .Q(\mem[170][10] ) );
  DFQD1 \mem_reg[170][9]  ( .D(n1942), .CP(clk), .Q(\mem[170][9] ) );
  DFQD1 \mem_reg[170][8]  ( .D(n1941), .CP(clk), .Q(\mem[170][8] ) );
  DFQD1 \mem_reg[170][7]  ( .D(n1940), .CP(clk), .Q(\mem[170][7] ) );
  DFQD1 \mem_reg[170][6]  ( .D(n1939), .CP(clk), .Q(\mem[170][6] ) );
  DFQD1 \mem_reg[170][5]  ( .D(n1938), .CP(clk), .Q(\mem[170][5] ) );
  DFQD1 \mem_reg[170][4]  ( .D(n1937), .CP(clk), .Q(\mem[170][4] ) );
  DFQD1 \mem_reg[170][3]  ( .D(n1936), .CP(clk), .Q(\mem[170][3] ) );
  DFQD1 \mem_reg[170][2]  ( .D(n1935), .CP(clk), .Q(\mem[170][2] ) );
  DFQD1 \mem_reg[170][1]  ( .D(n1934), .CP(clk), .Q(\mem[170][1] ) );
  DFQD1 \mem_reg[170][0]  ( .D(n1933), .CP(clk), .Q(\mem[170][0] ) );
  DFQD1 \mem_reg[171][15]  ( .D(n1932), .CP(clk), .Q(\mem[171][15] ) );
  DFQD1 \mem_reg[171][14]  ( .D(n1931), .CP(clk), .Q(\mem[171][14] ) );
  DFQD1 \mem_reg[171][13]  ( .D(n1930), .CP(clk), .Q(\mem[171][13] ) );
  DFQD1 \mem_reg[171][12]  ( .D(n1929), .CP(clk), .Q(\mem[171][12] ) );
  DFQD1 \mem_reg[171][11]  ( .D(n1928), .CP(clk), .Q(\mem[171][11] ) );
  DFQD1 \mem_reg[171][10]  ( .D(n1927), .CP(clk), .Q(\mem[171][10] ) );
  DFQD1 \mem_reg[171][9]  ( .D(n1926), .CP(clk), .Q(\mem[171][9] ) );
  DFQD1 \mem_reg[171][8]  ( .D(n1925), .CP(clk), .Q(\mem[171][8] ) );
  DFQD1 \mem_reg[171][7]  ( .D(n1924), .CP(clk), .Q(\mem[171][7] ) );
  DFQD1 \mem_reg[171][6]  ( .D(n1923), .CP(clk), .Q(\mem[171][6] ) );
  DFQD1 \mem_reg[171][5]  ( .D(n1922), .CP(clk), .Q(\mem[171][5] ) );
  DFQD1 \mem_reg[171][4]  ( .D(n1921), .CP(clk), .Q(\mem[171][4] ) );
  DFQD1 \mem_reg[171][3]  ( .D(n1920), .CP(clk), .Q(\mem[171][3] ) );
  DFQD1 \mem_reg[171][2]  ( .D(n1919), .CP(clk), .Q(\mem[171][2] ) );
  DFQD1 \mem_reg[171][1]  ( .D(n1918), .CP(clk), .Q(\mem[171][1] ) );
  DFQD1 \mem_reg[171][0]  ( .D(n1917), .CP(clk), .Q(\mem[171][0] ) );
  DFQD1 \mem_reg[172][15]  ( .D(n1916), .CP(clk), .Q(\mem[172][15] ) );
  DFQD1 \mem_reg[172][14]  ( .D(n1915), .CP(clk), .Q(\mem[172][14] ) );
  DFQD1 \mem_reg[172][13]  ( .D(n1914), .CP(clk), .Q(\mem[172][13] ) );
  DFQD1 \mem_reg[172][12]  ( .D(n1913), .CP(clk), .Q(\mem[172][12] ) );
  DFQD1 \mem_reg[172][11]  ( .D(n1912), .CP(clk), .Q(\mem[172][11] ) );
  DFQD1 \mem_reg[172][10]  ( .D(n1911), .CP(clk), .Q(\mem[172][10] ) );
  DFQD1 \mem_reg[172][9]  ( .D(n1910), .CP(clk), .Q(\mem[172][9] ) );
  DFQD1 \mem_reg[172][8]  ( .D(n1909), .CP(clk), .Q(\mem[172][8] ) );
  DFQD1 \mem_reg[172][7]  ( .D(n1908), .CP(clk), .Q(\mem[172][7] ) );
  DFQD1 \mem_reg[172][6]  ( .D(n1907), .CP(clk), .Q(\mem[172][6] ) );
  DFQD1 \mem_reg[172][5]  ( .D(n1906), .CP(clk), .Q(\mem[172][5] ) );
  DFQD1 \mem_reg[172][4]  ( .D(n1905), .CP(clk), .Q(\mem[172][4] ) );
  DFQD1 \mem_reg[172][3]  ( .D(n1904), .CP(clk), .Q(\mem[172][3] ) );
  DFQD1 \mem_reg[172][2]  ( .D(n1903), .CP(clk), .Q(\mem[172][2] ) );
  DFQD1 \mem_reg[172][1]  ( .D(n1902), .CP(clk), .Q(\mem[172][1] ) );
  DFQD1 \mem_reg[172][0]  ( .D(n1901), .CP(clk), .Q(\mem[172][0] ) );
  DFQD1 \mem_reg[173][15]  ( .D(n1900), .CP(clk), .Q(\mem[173][15] ) );
  DFQD1 \mem_reg[173][14]  ( .D(n1899), .CP(clk), .Q(\mem[173][14] ) );
  DFQD1 \mem_reg[173][13]  ( .D(n1898), .CP(clk), .Q(\mem[173][13] ) );
  DFQD1 \mem_reg[173][12]  ( .D(n1897), .CP(clk), .Q(\mem[173][12] ) );
  DFQD1 \mem_reg[173][11]  ( .D(n1896), .CP(clk), .Q(\mem[173][11] ) );
  DFQD1 \mem_reg[173][10]  ( .D(n1895), .CP(clk), .Q(\mem[173][10] ) );
  DFQD1 \mem_reg[173][9]  ( .D(n1894), .CP(clk), .Q(\mem[173][9] ) );
  DFQD1 \mem_reg[173][8]  ( .D(n1893), .CP(clk), .Q(\mem[173][8] ) );
  DFQD1 \mem_reg[173][7]  ( .D(n1892), .CP(clk), .Q(\mem[173][7] ) );
  DFQD1 \mem_reg[173][6]  ( .D(n1891), .CP(clk), .Q(\mem[173][6] ) );
  DFQD1 \mem_reg[173][5]  ( .D(n1890), .CP(clk), .Q(\mem[173][5] ) );
  DFQD1 \mem_reg[173][4]  ( .D(n1889), .CP(clk), .Q(\mem[173][4] ) );
  DFQD1 \mem_reg[173][3]  ( .D(n1888), .CP(clk), .Q(\mem[173][3] ) );
  DFQD1 \mem_reg[173][2]  ( .D(n1887), .CP(clk), .Q(\mem[173][2] ) );
  DFQD1 \mem_reg[173][1]  ( .D(n1886), .CP(clk), .Q(\mem[173][1] ) );
  DFQD1 \mem_reg[173][0]  ( .D(n1885), .CP(clk), .Q(\mem[173][0] ) );
  DFQD1 \mem_reg[174][15]  ( .D(n1884), .CP(clk), .Q(\mem[174][15] ) );
  DFQD1 \mem_reg[174][14]  ( .D(n1883), .CP(clk), .Q(\mem[174][14] ) );
  DFQD1 \mem_reg[174][13]  ( .D(n1882), .CP(clk), .Q(\mem[174][13] ) );
  DFQD1 \mem_reg[174][12]  ( .D(n1881), .CP(clk), .Q(\mem[174][12] ) );
  DFQD1 \mem_reg[174][11]  ( .D(n1880), .CP(clk), .Q(\mem[174][11] ) );
  DFQD1 \mem_reg[174][10]  ( .D(n1879), .CP(clk), .Q(\mem[174][10] ) );
  DFQD1 \mem_reg[174][9]  ( .D(n1878), .CP(clk), .Q(\mem[174][9] ) );
  DFQD1 \mem_reg[174][8]  ( .D(n1877), .CP(clk), .Q(\mem[174][8] ) );
  DFQD1 \mem_reg[174][7]  ( .D(n1876), .CP(clk), .Q(\mem[174][7] ) );
  DFQD1 \mem_reg[174][6]  ( .D(n1875), .CP(clk), .Q(\mem[174][6] ) );
  DFQD1 \mem_reg[174][5]  ( .D(n1874), .CP(clk), .Q(\mem[174][5] ) );
  DFQD1 \mem_reg[174][4]  ( .D(n1873), .CP(clk), .Q(\mem[174][4] ) );
  DFQD1 \mem_reg[174][3]  ( .D(n1872), .CP(clk), .Q(\mem[174][3] ) );
  DFQD1 \mem_reg[174][2]  ( .D(n1871), .CP(clk), .Q(\mem[174][2] ) );
  DFQD1 \mem_reg[174][1]  ( .D(n1870), .CP(clk), .Q(\mem[174][1] ) );
  DFQD1 \mem_reg[174][0]  ( .D(n1869), .CP(clk), .Q(\mem[174][0] ) );
  DFQD1 \mem_reg[175][15]  ( .D(n1868), .CP(clk), .Q(\mem[175][15] ) );
  DFQD1 \mem_reg[175][14]  ( .D(n1867), .CP(clk), .Q(\mem[175][14] ) );
  DFQD1 \mem_reg[175][13]  ( .D(n1866), .CP(clk), .Q(\mem[175][13] ) );
  DFQD1 \mem_reg[175][12]  ( .D(n1865), .CP(clk), .Q(\mem[175][12] ) );
  DFQD1 \mem_reg[175][11]  ( .D(n1864), .CP(clk), .Q(\mem[175][11] ) );
  DFQD1 \mem_reg[175][10]  ( .D(n1863), .CP(clk), .Q(\mem[175][10] ) );
  DFQD1 \mem_reg[175][9]  ( .D(n1862), .CP(clk), .Q(\mem[175][9] ) );
  DFQD1 \mem_reg[175][8]  ( .D(n1861), .CP(clk), .Q(\mem[175][8] ) );
  DFQD1 \mem_reg[175][7]  ( .D(n1860), .CP(clk), .Q(\mem[175][7] ) );
  DFQD1 \mem_reg[175][6]  ( .D(n1859), .CP(clk), .Q(\mem[175][6] ) );
  DFQD1 \mem_reg[175][5]  ( .D(n1858), .CP(clk), .Q(\mem[175][5] ) );
  DFQD1 \mem_reg[175][4]  ( .D(n1857), .CP(clk), .Q(\mem[175][4] ) );
  DFQD1 \mem_reg[175][3]  ( .D(n1856), .CP(clk), .Q(\mem[175][3] ) );
  DFQD1 \mem_reg[175][2]  ( .D(n1855), .CP(clk), .Q(\mem[175][2] ) );
  DFQD1 \mem_reg[175][1]  ( .D(n1854), .CP(clk), .Q(\mem[175][1] ) );
  DFQD1 \mem_reg[175][0]  ( .D(n1853), .CP(clk), .Q(\mem[175][0] ) );
  DFQD1 \mem_reg[176][15]  ( .D(n1852), .CP(clk), .Q(\mem[176][15] ) );
  DFQD1 \mem_reg[176][14]  ( .D(n1851), .CP(clk), .Q(\mem[176][14] ) );
  DFQD1 \mem_reg[176][13]  ( .D(n1850), .CP(clk), .Q(\mem[176][13] ) );
  DFQD1 \mem_reg[176][12]  ( .D(n1849), .CP(clk), .Q(\mem[176][12] ) );
  DFQD1 \mem_reg[176][11]  ( .D(n1848), .CP(clk), .Q(\mem[176][11] ) );
  DFQD1 \mem_reg[176][10]  ( .D(n1847), .CP(clk), .Q(\mem[176][10] ) );
  DFQD1 \mem_reg[176][9]  ( .D(n1846), .CP(clk), .Q(\mem[176][9] ) );
  DFQD1 \mem_reg[176][8]  ( .D(n1845), .CP(clk), .Q(\mem[176][8] ) );
  DFQD1 \mem_reg[176][7]  ( .D(n1844), .CP(clk), .Q(\mem[176][7] ) );
  DFQD1 \mem_reg[176][6]  ( .D(n1843), .CP(clk), .Q(\mem[176][6] ) );
  DFQD1 \mem_reg[176][5]  ( .D(n1842), .CP(clk), .Q(\mem[176][5] ) );
  DFQD1 \mem_reg[176][4]  ( .D(n1841), .CP(clk), .Q(\mem[176][4] ) );
  DFQD1 \mem_reg[176][3]  ( .D(n1840), .CP(clk), .Q(\mem[176][3] ) );
  DFQD1 \mem_reg[176][2]  ( .D(n1839), .CP(clk), .Q(\mem[176][2] ) );
  DFQD1 \mem_reg[176][1]  ( .D(n1838), .CP(clk), .Q(\mem[176][1] ) );
  DFQD1 \mem_reg[176][0]  ( .D(n1837), .CP(clk), .Q(\mem[176][0] ) );
  DFQD1 \mem_reg[177][15]  ( .D(n1836), .CP(clk), .Q(\mem[177][15] ) );
  DFQD1 \mem_reg[177][14]  ( .D(n1835), .CP(clk), .Q(\mem[177][14] ) );
  DFQD1 \mem_reg[177][13]  ( .D(n1834), .CP(clk), .Q(\mem[177][13] ) );
  DFQD1 \mem_reg[177][12]  ( .D(n1833), .CP(clk), .Q(\mem[177][12] ) );
  DFQD1 \mem_reg[177][11]  ( .D(n1832), .CP(clk), .Q(\mem[177][11] ) );
  DFQD1 \mem_reg[177][10]  ( .D(n1831), .CP(clk), .Q(\mem[177][10] ) );
  DFQD1 \mem_reg[177][9]  ( .D(n1830), .CP(clk), .Q(\mem[177][9] ) );
  DFQD1 \mem_reg[177][8]  ( .D(n1829), .CP(clk), .Q(\mem[177][8] ) );
  DFQD1 \mem_reg[177][7]  ( .D(n1828), .CP(clk), .Q(\mem[177][7] ) );
  DFQD1 \mem_reg[177][6]  ( .D(n1827), .CP(clk), .Q(\mem[177][6] ) );
  DFQD1 \mem_reg[177][5]  ( .D(n1826), .CP(clk), .Q(\mem[177][5] ) );
  DFQD1 \mem_reg[177][4]  ( .D(n1825), .CP(clk), .Q(\mem[177][4] ) );
  DFQD1 \mem_reg[177][3]  ( .D(n1824), .CP(clk), .Q(\mem[177][3] ) );
  DFQD1 \mem_reg[177][2]  ( .D(n1823), .CP(clk), .Q(\mem[177][2] ) );
  DFQD1 \mem_reg[177][1]  ( .D(n1822), .CP(clk), .Q(\mem[177][1] ) );
  DFQD1 \mem_reg[177][0]  ( .D(n1821), .CP(clk), .Q(\mem[177][0] ) );
  DFQD1 \mem_reg[178][15]  ( .D(n1820), .CP(clk), .Q(\mem[178][15] ) );
  DFQD1 \mem_reg[178][14]  ( .D(n1819), .CP(clk), .Q(\mem[178][14] ) );
  DFQD1 \mem_reg[178][13]  ( .D(n1818), .CP(clk), .Q(\mem[178][13] ) );
  DFQD1 \mem_reg[178][12]  ( .D(n1817), .CP(clk), .Q(\mem[178][12] ) );
  DFQD1 \mem_reg[178][11]  ( .D(n1816), .CP(clk), .Q(\mem[178][11] ) );
  DFQD1 \mem_reg[178][10]  ( .D(n1815), .CP(clk), .Q(\mem[178][10] ) );
  DFQD1 \mem_reg[178][9]  ( .D(n1814), .CP(clk), .Q(\mem[178][9] ) );
  DFQD1 \mem_reg[178][8]  ( .D(n1813), .CP(clk), .Q(\mem[178][8] ) );
  DFQD1 \mem_reg[178][7]  ( .D(n1812), .CP(clk), .Q(\mem[178][7] ) );
  DFQD1 \mem_reg[178][6]  ( .D(n1811), .CP(clk), .Q(\mem[178][6] ) );
  DFQD1 \mem_reg[178][5]  ( .D(n1810), .CP(clk), .Q(\mem[178][5] ) );
  DFQD1 \mem_reg[178][4]  ( .D(n1809), .CP(clk), .Q(\mem[178][4] ) );
  DFQD1 \mem_reg[178][3]  ( .D(n1808), .CP(clk), .Q(\mem[178][3] ) );
  DFQD1 \mem_reg[178][2]  ( .D(n1807), .CP(clk), .Q(\mem[178][2] ) );
  DFQD1 \mem_reg[178][1]  ( .D(n1806), .CP(clk), .Q(\mem[178][1] ) );
  DFQD1 \mem_reg[178][0]  ( .D(n1805), .CP(clk), .Q(\mem[178][0] ) );
  DFQD1 \mem_reg[179][15]  ( .D(n1804), .CP(clk), .Q(\mem[179][15] ) );
  DFQD1 \mem_reg[179][14]  ( .D(n1803), .CP(clk), .Q(\mem[179][14] ) );
  DFQD1 \mem_reg[179][13]  ( .D(n1802), .CP(clk), .Q(\mem[179][13] ) );
  DFQD1 \mem_reg[179][12]  ( .D(n1801), .CP(clk), .Q(\mem[179][12] ) );
  DFQD1 \mem_reg[179][11]  ( .D(n1800), .CP(clk), .Q(\mem[179][11] ) );
  DFQD1 \mem_reg[179][10]  ( .D(n1799), .CP(clk), .Q(\mem[179][10] ) );
  DFQD1 \mem_reg[179][9]  ( .D(n1798), .CP(clk), .Q(\mem[179][9] ) );
  DFQD1 \mem_reg[179][8]  ( .D(n1797), .CP(clk), .Q(\mem[179][8] ) );
  DFQD1 \mem_reg[179][7]  ( .D(n1796), .CP(clk), .Q(\mem[179][7] ) );
  DFQD1 \mem_reg[179][6]  ( .D(n1795), .CP(clk), .Q(\mem[179][6] ) );
  DFQD1 \mem_reg[179][5]  ( .D(n1794), .CP(clk), .Q(\mem[179][5] ) );
  DFQD1 \mem_reg[179][4]  ( .D(n1793), .CP(clk), .Q(\mem[179][4] ) );
  DFQD1 \mem_reg[179][3]  ( .D(n1792), .CP(clk), .Q(\mem[179][3] ) );
  DFQD1 \mem_reg[179][2]  ( .D(n1791), .CP(clk), .Q(\mem[179][2] ) );
  DFQD1 \mem_reg[179][1]  ( .D(n1790), .CP(clk), .Q(\mem[179][1] ) );
  DFQD1 \mem_reg[179][0]  ( .D(n1789), .CP(clk), .Q(\mem[179][0] ) );
  DFQD1 \mem_reg[180][15]  ( .D(n1788), .CP(clk), .Q(\mem[180][15] ) );
  DFQD1 \mem_reg[180][14]  ( .D(n1787), .CP(clk), .Q(\mem[180][14] ) );
  DFQD1 \mem_reg[180][13]  ( .D(n1786), .CP(clk), .Q(\mem[180][13] ) );
  DFQD1 \mem_reg[180][12]  ( .D(n1785), .CP(clk), .Q(\mem[180][12] ) );
  DFQD1 \mem_reg[180][11]  ( .D(n1784), .CP(clk), .Q(\mem[180][11] ) );
  DFQD1 \mem_reg[180][10]  ( .D(n1783), .CP(clk), .Q(\mem[180][10] ) );
  DFQD1 \mem_reg[180][9]  ( .D(n1782), .CP(clk), .Q(\mem[180][9] ) );
  DFQD1 \mem_reg[180][8]  ( .D(n1781), .CP(clk), .Q(\mem[180][8] ) );
  DFQD1 \mem_reg[180][7]  ( .D(n1780), .CP(clk), .Q(\mem[180][7] ) );
  DFQD1 \mem_reg[180][6]  ( .D(n1779), .CP(clk), .Q(\mem[180][6] ) );
  DFQD1 \mem_reg[180][5]  ( .D(n1778), .CP(clk), .Q(\mem[180][5] ) );
  DFQD1 \mem_reg[180][4]  ( .D(n1777), .CP(clk), .Q(\mem[180][4] ) );
  DFQD1 \mem_reg[180][3]  ( .D(n1776), .CP(clk), .Q(\mem[180][3] ) );
  DFQD1 \mem_reg[180][2]  ( .D(n1775), .CP(clk), .Q(\mem[180][2] ) );
  DFQD1 \mem_reg[180][1]  ( .D(n1774), .CP(clk), .Q(\mem[180][1] ) );
  DFQD1 \mem_reg[180][0]  ( .D(n1773), .CP(clk), .Q(\mem[180][0] ) );
  DFQD1 \mem_reg[181][15]  ( .D(n1772), .CP(clk), .Q(\mem[181][15] ) );
  DFQD1 \mem_reg[181][14]  ( .D(n1771), .CP(clk), .Q(\mem[181][14] ) );
  DFQD1 \mem_reg[181][13]  ( .D(n1770), .CP(clk), .Q(\mem[181][13] ) );
  DFQD1 \mem_reg[181][12]  ( .D(n1769), .CP(clk), .Q(\mem[181][12] ) );
  DFQD1 \mem_reg[181][11]  ( .D(n1768), .CP(clk), .Q(\mem[181][11] ) );
  DFQD1 \mem_reg[181][10]  ( .D(n1767), .CP(clk), .Q(\mem[181][10] ) );
  DFQD1 \mem_reg[181][9]  ( .D(n1766), .CP(clk), .Q(\mem[181][9] ) );
  DFQD1 \mem_reg[181][8]  ( .D(n1765), .CP(clk), .Q(\mem[181][8] ) );
  DFQD1 \mem_reg[181][7]  ( .D(n1764), .CP(clk), .Q(\mem[181][7] ) );
  DFQD1 \mem_reg[181][6]  ( .D(n1763), .CP(clk), .Q(\mem[181][6] ) );
  DFQD1 \mem_reg[181][5]  ( .D(n1762), .CP(clk), .Q(\mem[181][5] ) );
  DFQD1 \mem_reg[181][4]  ( .D(n1761), .CP(clk), .Q(\mem[181][4] ) );
  DFQD1 \mem_reg[181][3]  ( .D(n1760), .CP(clk), .Q(\mem[181][3] ) );
  DFQD1 \mem_reg[181][2]  ( .D(n1759), .CP(clk), .Q(\mem[181][2] ) );
  DFQD1 \mem_reg[181][1]  ( .D(n1758), .CP(clk), .Q(\mem[181][1] ) );
  DFQD1 \mem_reg[181][0]  ( .D(n1757), .CP(clk), .Q(\mem[181][0] ) );
  DFQD1 \mem_reg[182][15]  ( .D(n1756), .CP(clk), .Q(\mem[182][15] ) );
  DFQD1 \mem_reg[182][14]  ( .D(n1755), .CP(clk), .Q(\mem[182][14] ) );
  DFQD1 \mem_reg[182][13]  ( .D(n1754), .CP(clk), .Q(\mem[182][13] ) );
  DFQD1 \mem_reg[182][12]  ( .D(n1753), .CP(clk), .Q(\mem[182][12] ) );
  DFQD1 \mem_reg[182][11]  ( .D(n1752), .CP(clk), .Q(\mem[182][11] ) );
  DFQD1 \mem_reg[182][10]  ( .D(n1751), .CP(clk), .Q(\mem[182][10] ) );
  DFQD1 \mem_reg[182][9]  ( .D(n1750), .CP(clk), .Q(\mem[182][9] ) );
  DFQD1 \mem_reg[182][8]  ( .D(n1749), .CP(clk), .Q(\mem[182][8] ) );
  DFQD1 \mem_reg[182][7]  ( .D(n1748), .CP(clk), .Q(\mem[182][7] ) );
  DFQD1 \mem_reg[182][6]  ( .D(n1747), .CP(clk), .Q(\mem[182][6] ) );
  DFQD1 \mem_reg[182][5]  ( .D(n1746), .CP(clk), .Q(\mem[182][5] ) );
  DFQD1 \mem_reg[182][4]  ( .D(n1745), .CP(clk), .Q(\mem[182][4] ) );
  DFQD1 \mem_reg[182][3]  ( .D(n1744), .CP(clk), .Q(\mem[182][3] ) );
  DFQD1 \mem_reg[182][2]  ( .D(n1743), .CP(clk), .Q(\mem[182][2] ) );
  DFQD1 \mem_reg[182][1]  ( .D(n1742), .CP(clk), .Q(\mem[182][1] ) );
  DFQD1 \mem_reg[182][0]  ( .D(n1741), .CP(clk), .Q(\mem[182][0] ) );
  DFQD1 \mem_reg[183][15]  ( .D(n1740), .CP(clk), .Q(\mem[183][15] ) );
  DFQD1 \mem_reg[183][14]  ( .D(n1739), .CP(clk), .Q(\mem[183][14] ) );
  DFQD1 \mem_reg[183][13]  ( .D(n1738), .CP(clk), .Q(\mem[183][13] ) );
  DFQD1 \mem_reg[183][12]  ( .D(n1737), .CP(clk), .Q(\mem[183][12] ) );
  DFQD1 \mem_reg[183][11]  ( .D(n1736), .CP(clk), .Q(\mem[183][11] ) );
  DFQD1 \mem_reg[183][10]  ( .D(n1735), .CP(clk), .Q(\mem[183][10] ) );
  DFQD1 \mem_reg[183][9]  ( .D(n1734), .CP(clk), .Q(\mem[183][9] ) );
  DFQD1 \mem_reg[183][8]  ( .D(n1733), .CP(clk), .Q(\mem[183][8] ) );
  DFQD1 \mem_reg[183][7]  ( .D(n1732), .CP(clk), .Q(\mem[183][7] ) );
  DFQD1 \mem_reg[183][6]  ( .D(n1731), .CP(clk), .Q(\mem[183][6] ) );
  DFQD1 \mem_reg[183][5]  ( .D(n1730), .CP(clk), .Q(\mem[183][5] ) );
  DFQD1 \mem_reg[183][4]  ( .D(n1729), .CP(clk), .Q(\mem[183][4] ) );
  DFQD1 \mem_reg[183][3]  ( .D(n1728), .CP(clk), .Q(\mem[183][3] ) );
  DFQD1 \mem_reg[183][2]  ( .D(n1727), .CP(clk), .Q(\mem[183][2] ) );
  DFQD1 \mem_reg[183][1]  ( .D(n1726), .CP(clk), .Q(\mem[183][1] ) );
  DFQD1 \mem_reg[183][0]  ( .D(n1725), .CP(clk), .Q(\mem[183][0] ) );
  DFQD1 \mem_reg[184][15]  ( .D(n1724), .CP(clk), .Q(\mem[184][15] ) );
  DFQD1 \mem_reg[184][14]  ( .D(n1723), .CP(clk), .Q(\mem[184][14] ) );
  DFQD1 \mem_reg[184][13]  ( .D(n1722), .CP(clk), .Q(\mem[184][13] ) );
  DFQD1 \mem_reg[184][12]  ( .D(n1721), .CP(clk), .Q(\mem[184][12] ) );
  DFQD1 \mem_reg[184][11]  ( .D(n1720), .CP(clk), .Q(\mem[184][11] ) );
  DFQD1 \mem_reg[184][10]  ( .D(n1719), .CP(clk), .Q(\mem[184][10] ) );
  DFQD1 \mem_reg[184][9]  ( .D(n1718), .CP(clk), .Q(\mem[184][9] ) );
  DFQD1 \mem_reg[184][8]  ( .D(n1717), .CP(clk), .Q(\mem[184][8] ) );
  DFQD1 \mem_reg[184][7]  ( .D(n1716), .CP(clk), .Q(\mem[184][7] ) );
  DFQD1 \mem_reg[184][6]  ( .D(n1715), .CP(clk), .Q(\mem[184][6] ) );
  DFQD1 \mem_reg[184][5]  ( .D(n1714), .CP(clk), .Q(\mem[184][5] ) );
  DFQD1 \mem_reg[184][4]  ( .D(n1713), .CP(clk), .Q(\mem[184][4] ) );
  DFQD1 \mem_reg[184][3]  ( .D(n1712), .CP(clk), .Q(\mem[184][3] ) );
  DFQD1 \mem_reg[184][2]  ( .D(n1711), .CP(clk), .Q(\mem[184][2] ) );
  DFQD1 \mem_reg[184][1]  ( .D(n1710), .CP(clk), .Q(\mem[184][1] ) );
  DFQD1 \mem_reg[184][0]  ( .D(n1709), .CP(clk), .Q(\mem[184][0] ) );
  DFQD1 \mem_reg[185][15]  ( .D(n1708), .CP(clk), .Q(\mem[185][15] ) );
  DFQD1 \mem_reg[185][14]  ( .D(n1707), .CP(clk), .Q(\mem[185][14] ) );
  DFQD1 \mem_reg[185][13]  ( .D(n1706), .CP(clk), .Q(\mem[185][13] ) );
  DFQD1 \mem_reg[185][12]  ( .D(n1705), .CP(clk), .Q(\mem[185][12] ) );
  DFQD1 \mem_reg[185][11]  ( .D(n1704), .CP(clk), .Q(\mem[185][11] ) );
  DFQD1 \mem_reg[185][10]  ( .D(n1703), .CP(clk), .Q(\mem[185][10] ) );
  DFQD1 \mem_reg[185][9]  ( .D(n1702), .CP(clk), .Q(\mem[185][9] ) );
  DFQD1 \mem_reg[185][8]  ( .D(n1701), .CP(clk), .Q(\mem[185][8] ) );
  DFQD1 \mem_reg[185][7]  ( .D(n1700), .CP(clk), .Q(\mem[185][7] ) );
  DFQD1 \mem_reg[185][6]  ( .D(n1699), .CP(clk), .Q(\mem[185][6] ) );
  DFQD1 \mem_reg[185][5]  ( .D(n1698), .CP(clk), .Q(\mem[185][5] ) );
  DFQD1 \mem_reg[185][4]  ( .D(n1697), .CP(clk), .Q(\mem[185][4] ) );
  DFQD1 \mem_reg[185][3]  ( .D(n1696), .CP(clk), .Q(\mem[185][3] ) );
  DFQD1 \mem_reg[185][2]  ( .D(n1695), .CP(clk), .Q(\mem[185][2] ) );
  DFQD1 \mem_reg[185][1]  ( .D(n1694), .CP(clk), .Q(\mem[185][1] ) );
  DFQD1 \mem_reg[185][0]  ( .D(n1693), .CP(clk), .Q(\mem[185][0] ) );
  DFQD1 \mem_reg[186][15]  ( .D(n1692), .CP(clk), .Q(\mem[186][15] ) );
  DFQD1 \mem_reg[186][14]  ( .D(n1691), .CP(clk), .Q(\mem[186][14] ) );
  DFQD1 \mem_reg[186][13]  ( .D(n1690), .CP(clk), .Q(\mem[186][13] ) );
  DFQD1 \mem_reg[186][12]  ( .D(n1689), .CP(clk), .Q(\mem[186][12] ) );
  DFQD1 \mem_reg[186][11]  ( .D(n1688), .CP(clk), .Q(\mem[186][11] ) );
  DFQD1 \mem_reg[186][10]  ( .D(n1687), .CP(clk), .Q(\mem[186][10] ) );
  DFQD1 \mem_reg[186][9]  ( .D(n1686), .CP(clk), .Q(\mem[186][9] ) );
  DFQD1 \mem_reg[186][8]  ( .D(n1685), .CP(clk), .Q(\mem[186][8] ) );
  DFQD1 \mem_reg[186][7]  ( .D(n1684), .CP(clk), .Q(\mem[186][7] ) );
  DFQD1 \mem_reg[186][6]  ( .D(n1683), .CP(clk), .Q(\mem[186][6] ) );
  DFQD1 \mem_reg[186][5]  ( .D(n1682), .CP(clk), .Q(\mem[186][5] ) );
  DFQD1 \mem_reg[186][4]  ( .D(n1681), .CP(clk), .Q(\mem[186][4] ) );
  DFQD1 \mem_reg[186][3]  ( .D(n1680), .CP(clk), .Q(\mem[186][3] ) );
  DFQD1 \mem_reg[186][2]  ( .D(n1679), .CP(clk), .Q(\mem[186][2] ) );
  DFQD1 \mem_reg[186][1]  ( .D(n1678), .CP(clk), .Q(\mem[186][1] ) );
  DFQD1 \mem_reg[186][0]  ( .D(n1677), .CP(clk), .Q(\mem[186][0] ) );
  DFQD1 \mem_reg[187][15]  ( .D(n1676), .CP(clk), .Q(\mem[187][15] ) );
  DFQD1 \mem_reg[187][14]  ( .D(n1675), .CP(clk), .Q(\mem[187][14] ) );
  DFQD1 \mem_reg[187][13]  ( .D(n1674), .CP(clk), .Q(\mem[187][13] ) );
  DFQD1 \mem_reg[187][12]  ( .D(n1673), .CP(clk), .Q(\mem[187][12] ) );
  DFQD1 \mem_reg[187][11]  ( .D(n1672), .CP(clk), .Q(\mem[187][11] ) );
  DFQD1 \mem_reg[187][10]  ( .D(n1671), .CP(clk), .Q(\mem[187][10] ) );
  DFQD1 \mem_reg[187][9]  ( .D(n1670), .CP(clk), .Q(\mem[187][9] ) );
  DFQD1 \mem_reg[187][8]  ( .D(n1669), .CP(clk), .Q(\mem[187][8] ) );
  DFQD1 \mem_reg[187][7]  ( .D(n1668), .CP(clk), .Q(\mem[187][7] ) );
  DFQD1 \mem_reg[187][6]  ( .D(n1667), .CP(clk), .Q(\mem[187][6] ) );
  DFQD1 \mem_reg[187][5]  ( .D(n1666), .CP(clk), .Q(\mem[187][5] ) );
  DFQD1 \mem_reg[187][4]  ( .D(n1665), .CP(clk), .Q(\mem[187][4] ) );
  DFQD1 \mem_reg[187][3]  ( .D(n1664), .CP(clk), .Q(\mem[187][3] ) );
  DFQD1 \mem_reg[187][2]  ( .D(n1663), .CP(clk), .Q(\mem[187][2] ) );
  DFQD1 \mem_reg[187][1]  ( .D(n1662), .CP(clk), .Q(\mem[187][1] ) );
  DFQD1 \mem_reg[187][0]  ( .D(n1661), .CP(clk), .Q(\mem[187][0] ) );
  DFQD1 \mem_reg[188][15]  ( .D(n1660), .CP(clk), .Q(\mem[188][15] ) );
  DFQD1 \mem_reg[188][14]  ( .D(n1659), .CP(clk), .Q(\mem[188][14] ) );
  DFQD1 \mem_reg[188][13]  ( .D(n1658), .CP(clk), .Q(\mem[188][13] ) );
  DFQD1 \mem_reg[188][12]  ( .D(n1657), .CP(clk), .Q(\mem[188][12] ) );
  DFQD1 \mem_reg[188][11]  ( .D(n1656), .CP(clk), .Q(\mem[188][11] ) );
  DFQD1 \mem_reg[188][10]  ( .D(n1655), .CP(clk), .Q(\mem[188][10] ) );
  DFQD1 \mem_reg[188][9]  ( .D(n1654), .CP(clk), .Q(\mem[188][9] ) );
  DFQD1 \mem_reg[188][8]  ( .D(n1653), .CP(clk), .Q(\mem[188][8] ) );
  DFQD1 \mem_reg[188][7]  ( .D(n1652), .CP(clk), .Q(\mem[188][7] ) );
  DFQD1 \mem_reg[188][6]  ( .D(n1651), .CP(clk), .Q(\mem[188][6] ) );
  DFQD1 \mem_reg[188][5]  ( .D(n1650), .CP(clk), .Q(\mem[188][5] ) );
  DFQD1 \mem_reg[188][4]  ( .D(n1649), .CP(clk), .Q(\mem[188][4] ) );
  DFQD1 \mem_reg[188][3]  ( .D(n1648), .CP(clk), .Q(\mem[188][3] ) );
  DFQD1 \mem_reg[188][2]  ( .D(n1647), .CP(clk), .Q(\mem[188][2] ) );
  DFQD1 \mem_reg[188][1]  ( .D(n1646), .CP(clk), .Q(\mem[188][1] ) );
  DFQD1 \mem_reg[188][0]  ( .D(n1645), .CP(clk), .Q(\mem[188][0] ) );
  DFQD1 \mem_reg[189][15]  ( .D(n1644), .CP(clk), .Q(\mem[189][15] ) );
  DFQD1 \mem_reg[189][14]  ( .D(n1643), .CP(clk), .Q(\mem[189][14] ) );
  DFQD1 \mem_reg[189][13]  ( .D(n1642), .CP(clk), .Q(\mem[189][13] ) );
  DFQD1 \mem_reg[189][12]  ( .D(n1641), .CP(clk), .Q(\mem[189][12] ) );
  DFQD1 \mem_reg[189][11]  ( .D(n1640), .CP(clk), .Q(\mem[189][11] ) );
  DFQD1 \mem_reg[189][10]  ( .D(n1639), .CP(clk), .Q(\mem[189][10] ) );
  DFQD1 \mem_reg[189][9]  ( .D(n1638), .CP(clk), .Q(\mem[189][9] ) );
  DFQD1 \mem_reg[189][8]  ( .D(n1637), .CP(clk), .Q(\mem[189][8] ) );
  DFQD1 \mem_reg[189][7]  ( .D(n1636), .CP(clk), .Q(\mem[189][7] ) );
  DFQD1 \mem_reg[189][6]  ( .D(n1635), .CP(clk), .Q(\mem[189][6] ) );
  DFQD1 \mem_reg[189][5]  ( .D(n1634), .CP(clk), .Q(\mem[189][5] ) );
  DFQD1 \mem_reg[189][4]  ( .D(n1633), .CP(clk), .Q(\mem[189][4] ) );
  DFQD1 \mem_reg[189][3]  ( .D(n1632), .CP(clk), .Q(\mem[189][3] ) );
  DFQD1 \mem_reg[189][2]  ( .D(n1631), .CP(clk), .Q(\mem[189][2] ) );
  DFQD1 \mem_reg[189][1]  ( .D(n1630), .CP(clk), .Q(\mem[189][1] ) );
  DFQD1 \mem_reg[189][0]  ( .D(n1629), .CP(clk), .Q(\mem[189][0] ) );
  DFQD1 \mem_reg[190][15]  ( .D(n1628), .CP(clk), .Q(\mem[190][15] ) );
  DFQD1 \mem_reg[190][14]  ( .D(n1627), .CP(clk), .Q(\mem[190][14] ) );
  DFQD1 \mem_reg[190][13]  ( .D(n1626), .CP(clk), .Q(\mem[190][13] ) );
  DFQD1 \mem_reg[190][12]  ( .D(n1625), .CP(clk), .Q(\mem[190][12] ) );
  DFQD1 \mem_reg[190][11]  ( .D(n1624), .CP(clk), .Q(\mem[190][11] ) );
  DFQD1 \mem_reg[190][10]  ( .D(n1623), .CP(clk), .Q(\mem[190][10] ) );
  DFQD1 \mem_reg[190][9]  ( .D(n1622), .CP(clk), .Q(\mem[190][9] ) );
  DFQD1 \mem_reg[190][8]  ( .D(n1621), .CP(clk), .Q(\mem[190][8] ) );
  DFQD1 \mem_reg[190][7]  ( .D(n1620), .CP(clk), .Q(\mem[190][7] ) );
  DFQD1 \mem_reg[190][6]  ( .D(n1619), .CP(clk), .Q(\mem[190][6] ) );
  DFQD1 \mem_reg[190][5]  ( .D(n1618), .CP(clk), .Q(\mem[190][5] ) );
  DFQD1 \mem_reg[190][4]  ( .D(n1617), .CP(clk), .Q(\mem[190][4] ) );
  DFQD1 \mem_reg[190][3]  ( .D(n1616), .CP(clk), .Q(\mem[190][3] ) );
  DFQD1 \mem_reg[190][2]  ( .D(n1615), .CP(clk), .Q(\mem[190][2] ) );
  DFQD1 \mem_reg[190][1]  ( .D(n1614), .CP(clk), .Q(\mem[190][1] ) );
  DFQD1 \mem_reg[190][0]  ( .D(n1613), .CP(clk), .Q(\mem[190][0] ) );
  DFQD1 \mem_reg[191][15]  ( .D(n1612), .CP(clk), .Q(\mem[191][15] ) );
  DFQD1 \mem_reg[191][14]  ( .D(n1611), .CP(clk), .Q(\mem[191][14] ) );
  DFQD1 \mem_reg[191][13]  ( .D(n1610), .CP(clk), .Q(\mem[191][13] ) );
  DFQD1 \mem_reg[191][12]  ( .D(n1609), .CP(clk), .Q(\mem[191][12] ) );
  DFQD1 \mem_reg[191][11]  ( .D(n1608), .CP(clk), .Q(\mem[191][11] ) );
  DFQD1 \mem_reg[191][10]  ( .D(n1607), .CP(clk), .Q(\mem[191][10] ) );
  DFQD1 \mem_reg[191][9]  ( .D(n1606), .CP(clk), .Q(\mem[191][9] ) );
  DFQD1 \mem_reg[191][8]  ( .D(n1605), .CP(clk), .Q(\mem[191][8] ) );
  DFQD1 \mem_reg[191][7]  ( .D(n1604), .CP(clk), .Q(\mem[191][7] ) );
  DFQD1 \mem_reg[191][6]  ( .D(n1603), .CP(clk), .Q(\mem[191][6] ) );
  DFQD1 \mem_reg[191][5]  ( .D(n1602), .CP(clk), .Q(\mem[191][5] ) );
  DFQD1 \mem_reg[191][4]  ( .D(n1601), .CP(clk), .Q(\mem[191][4] ) );
  DFQD1 \mem_reg[191][3]  ( .D(n1600), .CP(clk), .Q(\mem[191][3] ) );
  DFQD1 \mem_reg[191][2]  ( .D(n1599), .CP(clk), .Q(\mem[191][2] ) );
  DFQD1 \mem_reg[191][1]  ( .D(n1598), .CP(clk), .Q(\mem[191][1] ) );
  DFQD1 \mem_reg[191][0]  ( .D(n1597), .CP(clk), .Q(\mem[191][0] ) );
  DFQD1 \mem_reg[192][15]  ( .D(n1596), .CP(clk), .Q(\mem[192][15] ) );
  DFQD1 \mem_reg[192][14]  ( .D(n1595), .CP(clk), .Q(\mem[192][14] ) );
  DFQD1 \mem_reg[192][13]  ( .D(n1594), .CP(clk), .Q(\mem[192][13] ) );
  DFQD1 \mem_reg[192][12]  ( .D(n1593), .CP(clk), .Q(\mem[192][12] ) );
  DFQD1 \mem_reg[192][11]  ( .D(n1592), .CP(clk), .Q(\mem[192][11] ) );
  DFQD1 \mem_reg[192][10]  ( .D(n1591), .CP(clk), .Q(\mem[192][10] ) );
  DFQD1 \mem_reg[192][9]  ( .D(n1590), .CP(clk), .Q(\mem[192][9] ) );
  DFQD1 \mem_reg[192][8]  ( .D(n1589), .CP(clk), .Q(\mem[192][8] ) );
  DFQD1 \mem_reg[192][7]  ( .D(n1588), .CP(clk), .Q(\mem[192][7] ) );
  DFQD1 \mem_reg[192][6]  ( .D(n1587), .CP(clk), .Q(\mem[192][6] ) );
  DFQD1 \mem_reg[192][5]  ( .D(n1586), .CP(clk), .Q(\mem[192][5] ) );
  DFQD1 \mem_reg[192][4]  ( .D(n1585), .CP(clk), .Q(\mem[192][4] ) );
  DFQD1 \mem_reg[192][3]  ( .D(n1584), .CP(clk), .Q(\mem[192][3] ) );
  DFQD1 \mem_reg[192][2]  ( .D(n1583), .CP(clk), .Q(\mem[192][2] ) );
  DFQD1 \mem_reg[192][1]  ( .D(n1582), .CP(clk), .Q(\mem[192][1] ) );
  DFQD1 \mem_reg[192][0]  ( .D(n1581), .CP(clk), .Q(\mem[192][0] ) );
  DFQD1 \mem_reg[193][15]  ( .D(n1580), .CP(clk), .Q(\mem[193][15] ) );
  DFQD1 \mem_reg[193][14]  ( .D(n1579), .CP(clk), .Q(\mem[193][14] ) );
  DFQD1 \mem_reg[193][13]  ( .D(n1578), .CP(clk), .Q(\mem[193][13] ) );
  DFQD1 \mem_reg[193][12]  ( .D(n1577), .CP(clk), .Q(\mem[193][12] ) );
  DFQD1 \mem_reg[193][11]  ( .D(n1576), .CP(clk), .Q(\mem[193][11] ) );
  DFQD1 \mem_reg[193][10]  ( .D(n1575), .CP(clk), .Q(\mem[193][10] ) );
  DFQD1 \mem_reg[193][9]  ( .D(n1574), .CP(clk), .Q(\mem[193][9] ) );
  DFQD1 \mem_reg[193][8]  ( .D(n1573), .CP(clk), .Q(\mem[193][8] ) );
  DFQD1 \mem_reg[193][7]  ( .D(n1572), .CP(clk), .Q(\mem[193][7] ) );
  DFQD1 \mem_reg[193][6]  ( .D(n1571), .CP(clk), .Q(\mem[193][6] ) );
  DFQD1 \mem_reg[193][5]  ( .D(n1570), .CP(clk), .Q(\mem[193][5] ) );
  DFQD1 \mem_reg[193][4]  ( .D(n1569), .CP(clk), .Q(\mem[193][4] ) );
  DFQD1 \mem_reg[193][3]  ( .D(n1568), .CP(clk), .Q(\mem[193][3] ) );
  DFQD1 \mem_reg[193][2]  ( .D(n1567), .CP(clk), .Q(\mem[193][2] ) );
  DFQD1 \mem_reg[193][1]  ( .D(n1566), .CP(clk), .Q(\mem[193][1] ) );
  DFQD1 \mem_reg[193][0]  ( .D(n1565), .CP(clk), .Q(\mem[193][0] ) );
  DFQD1 \mem_reg[194][15]  ( .D(n1564), .CP(clk), .Q(\mem[194][15] ) );
  DFQD1 \mem_reg[194][14]  ( .D(n1563), .CP(clk), .Q(\mem[194][14] ) );
  DFQD1 \mem_reg[194][13]  ( .D(n1562), .CP(clk), .Q(\mem[194][13] ) );
  DFQD1 \mem_reg[194][12]  ( .D(n1561), .CP(clk), .Q(\mem[194][12] ) );
  DFQD1 \mem_reg[194][11]  ( .D(n1560), .CP(clk), .Q(\mem[194][11] ) );
  DFQD1 \mem_reg[194][10]  ( .D(n1559), .CP(clk), .Q(\mem[194][10] ) );
  DFQD1 \mem_reg[194][9]  ( .D(n1558), .CP(clk), .Q(\mem[194][9] ) );
  DFQD1 \mem_reg[194][8]  ( .D(n1557), .CP(clk), .Q(\mem[194][8] ) );
  DFQD1 \mem_reg[194][7]  ( .D(n1556), .CP(clk), .Q(\mem[194][7] ) );
  DFQD1 \mem_reg[194][6]  ( .D(n1555), .CP(clk), .Q(\mem[194][6] ) );
  DFQD1 \mem_reg[194][5]  ( .D(n1554), .CP(clk), .Q(\mem[194][5] ) );
  DFQD1 \mem_reg[194][4]  ( .D(n1553), .CP(clk), .Q(\mem[194][4] ) );
  DFQD1 \mem_reg[194][3]  ( .D(n1552), .CP(clk), .Q(\mem[194][3] ) );
  DFQD1 \mem_reg[194][2]  ( .D(n1551), .CP(clk), .Q(\mem[194][2] ) );
  DFQD1 \mem_reg[194][1]  ( .D(n1550), .CP(clk), .Q(\mem[194][1] ) );
  DFQD1 \mem_reg[194][0]  ( .D(n1549), .CP(clk), .Q(\mem[194][0] ) );
  DFQD1 \mem_reg[195][15]  ( .D(n1548), .CP(clk), .Q(\mem[195][15] ) );
  DFQD1 \mem_reg[195][14]  ( .D(n1547), .CP(clk), .Q(\mem[195][14] ) );
  DFQD1 \mem_reg[195][13]  ( .D(n1546), .CP(clk), .Q(\mem[195][13] ) );
  DFQD1 \mem_reg[195][12]  ( .D(n1545), .CP(clk), .Q(\mem[195][12] ) );
  DFQD1 \mem_reg[195][11]  ( .D(n1544), .CP(clk), .Q(\mem[195][11] ) );
  DFQD1 \mem_reg[195][10]  ( .D(n1543), .CP(clk), .Q(\mem[195][10] ) );
  DFQD1 \mem_reg[195][9]  ( .D(n1542), .CP(clk), .Q(\mem[195][9] ) );
  DFQD1 \mem_reg[195][8]  ( .D(n1541), .CP(clk), .Q(\mem[195][8] ) );
  DFQD1 \mem_reg[195][7]  ( .D(n1540), .CP(clk), .Q(\mem[195][7] ) );
  DFQD1 \mem_reg[195][6]  ( .D(n1539), .CP(clk), .Q(\mem[195][6] ) );
  DFQD1 \mem_reg[195][5]  ( .D(n1538), .CP(clk), .Q(\mem[195][5] ) );
  DFQD1 \mem_reg[195][4]  ( .D(n1537), .CP(clk), .Q(\mem[195][4] ) );
  DFQD1 \mem_reg[195][3]  ( .D(n1536), .CP(clk), .Q(\mem[195][3] ) );
  DFQD1 \mem_reg[195][2]  ( .D(n1535), .CP(clk), .Q(\mem[195][2] ) );
  DFQD1 \mem_reg[195][1]  ( .D(n1534), .CP(clk), .Q(\mem[195][1] ) );
  DFQD1 \mem_reg[195][0]  ( .D(n1533), .CP(clk), .Q(\mem[195][0] ) );
  DFQD1 \mem_reg[196][15]  ( .D(n1532), .CP(clk), .Q(\mem[196][15] ) );
  DFQD1 \mem_reg[196][14]  ( .D(n1531), .CP(clk), .Q(\mem[196][14] ) );
  DFQD1 \mem_reg[196][13]  ( .D(n1530), .CP(clk), .Q(\mem[196][13] ) );
  DFQD1 \mem_reg[196][12]  ( .D(n1529), .CP(clk), .Q(\mem[196][12] ) );
  DFQD1 \mem_reg[196][11]  ( .D(n1528), .CP(clk), .Q(\mem[196][11] ) );
  DFQD1 \mem_reg[196][10]  ( .D(n1527), .CP(clk), .Q(\mem[196][10] ) );
  DFQD1 \mem_reg[196][9]  ( .D(n1526), .CP(clk), .Q(\mem[196][9] ) );
  DFQD1 \mem_reg[196][8]  ( .D(n1525), .CP(clk), .Q(\mem[196][8] ) );
  DFQD1 \mem_reg[196][7]  ( .D(n1524), .CP(clk), .Q(\mem[196][7] ) );
  DFQD1 \mem_reg[196][6]  ( .D(n1523), .CP(clk), .Q(\mem[196][6] ) );
  DFQD1 \mem_reg[196][5]  ( .D(n1522), .CP(clk), .Q(\mem[196][5] ) );
  DFQD1 \mem_reg[196][4]  ( .D(n1521), .CP(clk), .Q(\mem[196][4] ) );
  DFQD1 \mem_reg[196][3]  ( .D(n1520), .CP(clk), .Q(\mem[196][3] ) );
  DFQD1 \mem_reg[196][2]  ( .D(n1519), .CP(clk), .Q(\mem[196][2] ) );
  DFQD1 \mem_reg[196][1]  ( .D(n1518), .CP(clk), .Q(\mem[196][1] ) );
  DFQD1 \mem_reg[196][0]  ( .D(n1517), .CP(clk), .Q(\mem[196][0] ) );
  DFQD1 \mem_reg[197][15]  ( .D(n1516), .CP(clk), .Q(\mem[197][15] ) );
  DFQD1 \mem_reg[197][14]  ( .D(n1515), .CP(clk), .Q(\mem[197][14] ) );
  DFQD1 \mem_reg[197][13]  ( .D(n1514), .CP(clk), .Q(\mem[197][13] ) );
  DFQD1 \mem_reg[197][12]  ( .D(n1513), .CP(clk), .Q(\mem[197][12] ) );
  DFQD1 \mem_reg[197][11]  ( .D(n1512), .CP(clk), .Q(\mem[197][11] ) );
  DFQD1 \mem_reg[197][10]  ( .D(n1511), .CP(clk), .Q(\mem[197][10] ) );
  DFQD1 \mem_reg[197][9]  ( .D(n1510), .CP(clk), .Q(\mem[197][9] ) );
  DFQD1 \mem_reg[197][8]  ( .D(n1509), .CP(clk), .Q(\mem[197][8] ) );
  DFQD1 \mem_reg[197][7]  ( .D(n1508), .CP(clk), .Q(\mem[197][7] ) );
  DFQD1 \mem_reg[197][6]  ( .D(n1507), .CP(clk), .Q(\mem[197][6] ) );
  DFQD1 \mem_reg[197][5]  ( .D(n1506), .CP(clk), .Q(\mem[197][5] ) );
  DFQD1 \mem_reg[197][4]  ( .D(n1505), .CP(clk), .Q(\mem[197][4] ) );
  DFQD1 \mem_reg[197][3]  ( .D(n1504), .CP(clk), .Q(\mem[197][3] ) );
  DFQD1 \mem_reg[197][2]  ( .D(n1503), .CP(clk), .Q(\mem[197][2] ) );
  DFQD1 \mem_reg[197][1]  ( .D(n1502), .CP(clk), .Q(\mem[197][1] ) );
  DFQD1 \mem_reg[197][0]  ( .D(n1501), .CP(clk), .Q(\mem[197][0] ) );
  DFQD1 \mem_reg[198][15]  ( .D(n1500), .CP(clk), .Q(\mem[198][15] ) );
  DFQD1 \mem_reg[198][14]  ( .D(n1499), .CP(clk), .Q(\mem[198][14] ) );
  DFQD1 \mem_reg[198][13]  ( .D(n1498), .CP(clk), .Q(\mem[198][13] ) );
  DFQD1 \mem_reg[198][12]  ( .D(n1497), .CP(clk), .Q(\mem[198][12] ) );
  DFQD1 \mem_reg[198][11]  ( .D(n1496), .CP(clk), .Q(\mem[198][11] ) );
  DFQD1 \mem_reg[198][10]  ( .D(n1495), .CP(clk), .Q(\mem[198][10] ) );
  DFQD1 \mem_reg[198][9]  ( .D(n1494), .CP(clk), .Q(\mem[198][9] ) );
  DFQD1 \mem_reg[198][8]  ( .D(n1493), .CP(clk), .Q(\mem[198][8] ) );
  DFQD1 \mem_reg[198][7]  ( .D(n1492), .CP(clk), .Q(\mem[198][7] ) );
  DFQD1 \mem_reg[198][6]  ( .D(n1491), .CP(clk), .Q(\mem[198][6] ) );
  DFQD1 \mem_reg[198][5]  ( .D(n1490), .CP(clk), .Q(\mem[198][5] ) );
  DFQD1 \mem_reg[198][4]  ( .D(n1489), .CP(clk), .Q(\mem[198][4] ) );
  DFQD1 \mem_reg[198][3]  ( .D(n1488), .CP(clk), .Q(\mem[198][3] ) );
  DFQD1 \mem_reg[198][2]  ( .D(n1487), .CP(clk), .Q(\mem[198][2] ) );
  DFQD1 \mem_reg[198][1]  ( .D(n1486), .CP(clk), .Q(\mem[198][1] ) );
  DFQD1 \mem_reg[198][0]  ( .D(n1485), .CP(clk), .Q(\mem[198][0] ) );
  DFQD1 \mem_reg[199][15]  ( .D(n1484), .CP(clk), .Q(\mem[199][15] ) );
  DFQD1 \mem_reg[199][14]  ( .D(n1483), .CP(clk), .Q(\mem[199][14] ) );
  DFQD1 \mem_reg[199][13]  ( .D(n1482), .CP(clk), .Q(\mem[199][13] ) );
  DFQD1 \mem_reg[199][12]  ( .D(n1481), .CP(clk), .Q(\mem[199][12] ) );
  DFQD1 \mem_reg[199][11]  ( .D(n1480), .CP(clk), .Q(\mem[199][11] ) );
  DFQD1 \mem_reg[199][10]  ( .D(n1479), .CP(clk), .Q(\mem[199][10] ) );
  DFQD1 \mem_reg[199][9]  ( .D(n1478), .CP(clk), .Q(\mem[199][9] ) );
  DFQD1 \mem_reg[199][8]  ( .D(n1477), .CP(clk), .Q(\mem[199][8] ) );
  DFQD1 \mem_reg[199][7]  ( .D(n1476), .CP(clk), .Q(\mem[199][7] ) );
  DFQD1 \mem_reg[199][6]  ( .D(n1475), .CP(clk), .Q(\mem[199][6] ) );
  DFQD1 \mem_reg[199][5]  ( .D(n1474), .CP(clk), .Q(\mem[199][5] ) );
  DFQD1 \mem_reg[199][4]  ( .D(n1473), .CP(clk), .Q(\mem[199][4] ) );
  DFQD1 \mem_reg[199][3]  ( .D(n1472), .CP(clk), .Q(\mem[199][3] ) );
  DFQD1 \mem_reg[199][2]  ( .D(n1471), .CP(clk), .Q(\mem[199][2] ) );
  DFQD1 \mem_reg[199][1]  ( .D(n1470), .CP(clk), .Q(\mem[199][1] ) );
  DFQD1 \mem_reg[199][0]  ( .D(n1469), .CP(clk), .Q(\mem[199][0] ) );
  DFQD1 \mem_reg[200][15]  ( .D(n1468), .CP(clk), .Q(\mem[200][15] ) );
  DFQD1 \mem_reg[200][14]  ( .D(n1467), .CP(clk), .Q(\mem[200][14] ) );
  DFQD1 \mem_reg[200][13]  ( .D(n1466), .CP(clk), .Q(\mem[200][13] ) );
  DFQD1 \mem_reg[200][12]  ( .D(n1465), .CP(clk), .Q(\mem[200][12] ) );
  DFQD1 \mem_reg[200][11]  ( .D(n1464), .CP(clk), .Q(\mem[200][11] ) );
  DFQD1 \mem_reg[200][10]  ( .D(n1463), .CP(clk), .Q(\mem[200][10] ) );
  DFQD1 \mem_reg[200][9]  ( .D(n1462), .CP(clk), .Q(\mem[200][9] ) );
  DFQD1 \mem_reg[200][8]  ( .D(n1461), .CP(clk), .Q(\mem[200][8] ) );
  DFQD1 \mem_reg[200][7]  ( .D(n1460), .CP(clk), .Q(\mem[200][7] ) );
  DFQD1 \mem_reg[200][6]  ( .D(n1459), .CP(clk), .Q(\mem[200][6] ) );
  DFQD1 \mem_reg[200][5]  ( .D(n1458), .CP(clk), .Q(\mem[200][5] ) );
  DFQD1 \mem_reg[200][4]  ( .D(n1457), .CP(clk), .Q(\mem[200][4] ) );
  DFQD1 \mem_reg[200][3]  ( .D(n1456), .CP(clk), .Q(\mem[200][3] ) );
  DFQD1 \mem_reg[200][2]  ( .D(n1455), .CP(clk), .Q(\mem[200][2] ) );
  DFQD1 \mem_reg[200][1]  ( .D(n1454), .CP(clk), .Q(\mem[200][1] ) );
  DFQD1 \mem_reg[200][0]  ( .D(n1453), .CP(clk), .Q(\mem[200][0] ) );
  DFQD1 \mem_reg[201][15]  ( .D(n1452), .CP(clk), .Q(\mem[201][15] ) );
  DFQD1 \mem_reg[201][14]  ( .D(n1451), .CP(clk), .Q(\mem[201][14] ) );
  DFQD1 \mem_reg[201][13]  ( .D(n1450), .CP(clk), .Q(\mem[201][13] ) );
  DFQD1 \mem_reg[201][12]  ( .D(n1449), .CP(clk), .Q(\mem[201][12] ) );
  DFQD1 \mem_reg[201][11]  ( .D(n1448), .CP(clk), .Q(\mem[201][11] ) );
  DFQD1 \mem_reg[201][10]  ( .D(n1447), .CP(clk), .Q(\mem[201][10] ) );
  DFQD1 \mem_reg[201][9]  ( .D(n1446), .CP(clk), .Q(\mem[201][9] ) );
  DFQD1 \mem_reg[201][8]  ( .D(n1445), .CP(clk), .Q(\mem[201][8] ) );
  DFQD1 \mem_reg[201][7]  ( .D(n1444), .CP(clk), .Q(\mem[201][7] ) );
  DFQD1 \mem_reg[201][6]  ( .D(n1443), .CP(clk), .Q(\mem[201][6] ) );
  DFQD1 \mem_reg[201][5]  ( .D(n1442), .CP(clk), .Q(\mem[201][5] ) );
  DFQD1 \mem_reg[201][4]  ( .D(n1441), .CP(clk), .Q(\mem[201][4] ) );
  DFQD1 \mem_reg[201][3]  ( .D(n1440), .CP(clk), .Q(\mem[201][3] ) );
  DFQD1 \mem_reg[201][2]  ( .D(n1439), .CP(clk), .Q(\mem[201][2] ) );
  DFQD1 \mem_reg[201][1]  ( .D(n1438), .CP(clk), .Q(\mem[201][1] ) );
  DFQD1 \mem_reg[201][0]  ( .D(n1437), .CP(clk), .Q(\mem[201][0] ) );
  DFQD1 \mem_reg[202][15]  ( .D(n1436), .CP(clk), .Q(\mem[202][15] ) );
  DFQD1 \mem_reg[202][14]  ( .D(n1435), .CP(clk), .Q(\mem[202][14] ) );
  DFQD1 \mem_reg[202][13]  ( .D(n1434), .CP(clk), .Q(\mem[202][13] ) );
  DFQD1 \mem_reg[202][12]  ( .D(n1433), .CP(clk), .Q(\mem[202][12] ) );
  DFQD1 \mem_reg[202][11]  ( .D(n1432), .CP(clk), .Q(\mem[202][11] ) );
  DFQD1 \mem_reg[202][10]  ( .D(n1431), .CP(clk), .Q(\mem[202][10] ) );
  DFQD1 \mem_reg[202][9]  ( .D(n1430), .CP(clk), .Q(\mem[202][9] ) );
  DFQD1 \mem_reg[202][8]  ( .D(n1429), .CP(clk), .Q(\mem[202][8] ) );
  DFQD1 \mem_reg[202][7]  ( .D(n1428), .CP(clk), .Q(\mem[202][7] ) );
  DFQD1 \mem_reg[202][6]  ( .D(n1427), .CP(clk), .Q(\mem[202][6] ) );
  DFQD1 \mem_reg[202][5]  ( .D(n1426), .CP(clk), .Q(\mem[202][5] ) );
  DFQD1 \mem_reg[202][4]  ( .D(n1425), .CP(clk), .Q(\mem[202][4] ) );
  DFQD1 \mem_reg[202][3]  ( .D(n1424), .CP(clk), .Q(\mem[202][3] ) );
  DFQD1 \mem_reg[202][2]  ( .D(n1423), .CP(clk), .Q(\mem[202][2] ) );
  DFQD1 \mem_reg[202][1]  ( .D(n1422), .CP(clk), .Q(\mem[202][1] ) );
  DFQD1 \mem_reg[202][0]  ( .D(n1421), .CP(clk), .Q(\mem[202][0] ) );
  DFQD1 \mem_reg[203][15]  ( .D(n1420), .CP(clk), .Q(\mem[203][15] ) );
  DFQD1 \mem_reg[203][14]  ( .D(n1419), .CP(clk), .Q(\mem[203][14] ) );
  DFQD1 \mem_reg[203][13]  ( .D(n1418), .CP(clk), .Q(\mem[203][13] ) );
  DFQD1 \mem_reg[203][12]  ( .D(n1417), .CP(clk), .Q(\mem[203][12] ) );
  DFQD1 \mem_reg[203][11]  ( .D(n1416), .CP(clk), .Q(\mem[203][11] ) );
  DFQD1 \mem_reg[203][10]  ( .D(n1415), .CP(clk), .Q(\mem[203][10] ) );
  DFQD1 \mem_reg[203][9]  ( .D(n1414), .CP(clk), .Q(\mem[203][9] ) );
  DFQD1 \mem_reg[203][8]  ( .D(n1413), .CP(clk), .Q(\mem[203][8] ) );
  DFQD1 \mem_reg[203][7]  ( .D(n1412), .CP(clk), .Q(\mem[203][7] ) );
  DFQD1 \mem_reg[203][6]  ( .D(n1411), .CP(clk), .Q(\mem[203][6] ) );
  DFQD1 \mem_reg[203][5]  ( .D(n1410), .CP(clk), .Q(\mem[203][5] ) );
  DFQD1 \mem_reg[203][4]  ( .D(n1409), .CP(clk), .Q(\mem[203][4] ) );
  DFQD1 \mem_reg[203][3]  ( .D(n1408), .CP(clk), .Q(\mem[203][3] ) );
  DFQD1 \mem_reg[203][2]  ( .D(n1407), .CP(clk), .Q(\mem[203][2] ) );
  DFQD1 \mem_reg[203][1]  ( .D(n1406), .CP(clk), .Q(\mem[203][1] ) );
  DFQD1 \mem_reg[203][0]  ( .D(n1405), .CP(clk), .Q(\mem[203][0] ) );
  DFQD1 \mem_reg[204][15]  ( .D(n1404), .CP(clk), .Q(\mem[204][15] ) );
  DFQD1 \mem_reg[204][14]  ( .D(n1403), .CP(clk), .Q(\mem[204][14] ) );
  DFQD1 \mem_reg[204][13]  ( .D(n1402), .CP(clk), .Q(\mem[204][13] ) );
  DFQD1 \mem_reg[204][12]  ( .D(n1401), .CP(clk), .Q(\mem[204][12] ) );
  DFQD1 \mem_reg[204][11]  ( .D(n1400), .CP(clk), .Q(\mem[204][11] ) );
  DFQD1 \mem_reg[204][10]  ( .D(n1399), .CP(clk), .Q(\mem[204][10] ) );
  DFQD1 \mem_reg[204][9]  ( .D(n1398), .CP(clk), .Q(\mem[204][9] ) );
  DFQD1 \mem_reg[204][8]  ( .D(n1397), .CP(clk), .Q(\mem[204][8] ) );
  DFQD1 \mem_reg[204][7]  ( .D(n1396), .CP(clk), .Q(\mem[204][7] ) );
  DFQD1 \mem_reg[204][6]  ( .D(n1395), .CP(clk), .Q(\mem[204][6] ) );
  DFQD1 \mem_reg[204][5]  ( .D(n1394), .CP(clk), .Q(\mem[204][5] ) );
  DFQD1 \mem_reg[204][4]  ( .D(n1393), .CP(clk), .Q(\mem[204][4] ) );
  DFQD1 \mem_reg[204][3]  ( .D(n1392), .CP(clk), .Q(\mem[204][3] ) );
  DFQD1 \mem_reg[204][2]  ( .D(n1391), .CP(clk), .Q(\mem[204][2] ) );
  DFQD1 \mem_reg[204][1]  ( .D(n1390), .CP(clk), .Q(\mem[204][1] ) );
  DFQD1 \mem_reg[204][0]  ( .D(n1389), .CP(clk), .Q(\mem[204][0] ) );
  DFQD1 \mem_reg[205][15]  ( .D(n1388), .CP(clk), .Q(\mem[205][15] ) );
  DFQD1 \mem_reg[205][14]  ( .D(n1387), .CP(clk), .Q(\mem[205][14] ) );
  DFQD1 \mem_reg[205][13]  ( .D(n1386), .CP(clk), .Q(\mem[205][13] ) );
  DFQD1 \mem_reg[205][12]  ( .D(n1385), .CP(clk), .Q(\mem[205][12] ) );
  DFQD1 \mem_reg[205][11]  ( .D(n1384), .CP(clk), .Q(\mem[205][11] ) );
  DFQD1 \mem_reg[205][10]  ( .D(n1383), .CP(clk), .Q(\mem[205][10] ) );
  DFQD1 \mem_reg[205][9]  ( .D(n1382), .CP(clk), .Q(\mem[205][9] ) );
  DFQD1 \mem_reg[205][8]  ( .D(n1381), .CP(clk), .Q(\mem[205][8] ) );
  DFQD1 \mem_reg[205][7]  ( .D(n1380), .CP(clk), .Q(\mem[205][7] ) );
  DFQD1 \mem_reg[205][6]  ( .D(n1379), .CP(clk), .Q(\mem[205][6] ) );
  DFQD1 \mem_reg[205][5]  ( .D(n1378), .CP(clk), .Q(\mem[205][5] ) );
  DFQD1 \mem_reg[205][4]  ( .D(n1377), .CP(clk), .Q(\mem[205][4] ) );
  DFQD1 \mem_reg[205][3]  ( .D(n1376), .CP(clk), .Q(\mem[205][3] ) );
  DFQD1 \mem_reg[205][2]  ( .D(n1375), .CP(clk), .Q(\mem[205][2] ) );
  DFQD1 \mem_reg[205][1]  ( .D(n1374), .CP(clk), .Q(\mem[205][1] ) );
  DFQD1 \mem_reg[205][0]  ( .D(n1373), .CP(clk), .Q(\mem[205][0] ) );
  DFQD1 \mem_reg[206][15]  ( .D(n1372), .CP(clk), .Q(\mem[206][15] ) );
  DFQD1 \mem_reg[206][14]  ( .D(n1371), .CP(clk), .Q(\mem[206][14] ) );
  DFQD1 \mem_reg[206][13]  ( .D(n1370), .CP(clk), .Q(\mem[206][13] ) );
  DFQD1 \mem_reg[206][12]  ( .D(n1369), .CP(clk), .Q(\mem[206][12] ) );
  DFQD1 \mem_reg[206][11]  ( .D(n1368), .CP(clk), .Q(\mem[206][11] ) );
  DFQD1 \mem_reg[206][10]  ( .D(n1367), .CP(clk), .Q(\mem[206][10] ) );
  DFQD1 \mem_reg[206][9]  ( .D(n1366), .CP(clk), .Q(\mem[206][9] ) );
  DFQD1 \mem_reg[206][8]  ( .D(n1365), .CP(clk), .Q(\mem[206][8] ) );
  DFQD1 \mem_reg[206][7]  ( .D(n1364), .CP(clk), .Q(\mem[206][7] ) );
  DFQD1 \mem_reg[206][6]  ( .D(n1363), .CP(clk), .Q(\mem[206][6] ) );
  DFQD1 \mem_reg[206][5]  ( .D(n1362), .CP(clk), .Q(\mem[206][5] ) );
  DFQD1 \mem_reg[206][4]  ( .D(n1361), .CP(clk), .Q(\mem[206][4] ) );
  DFQD1 \mem_reg[206][3]  ( .D(n1360), .CP(clk), .Q(\mem[206][3] ) );
  DFQD1 \mem_reg[206][2]  ( .D(n1359), .CP(clk), .Q(\mem[206][2] ) );
  DFQD1 \mem_reg[206][1]  ( .D(n1358), .CP(clk), .Q(\mem[206][1] ) );
  DFQD1 \mem_reg[206][0]  ( .D(n1357), .CP(clk), .Q(\mem[206][0] ) );
  DFQD1 \mem_reg[207][15]  ( .D(n1356), .CP(clk), .Q(\mem[207][15] ) );
  DFQD1 \mem_reg[207][14]  ( .D(n1355), .CP(clk), .Q(\mem[207][14] ) );
  DFQD1 \mem_reg[207][13]  ( .D(n1354), .CP(clk), .Q(\mem[207][13] ) );
  DFQD1 \mem_reg[207][12]  ( .D(n1353), .CP(clk), .Q(\mem[207][12] ) );
  DFQD1 \mem_reg[207][11]  ( .D(n1352), .CP(clk), .Q(\mem[207][11] ) );
  DFQD1 \mem_reg[207][10]  ( .D(n1351), .CP(clk), .Q(\mem[207][10] ) );
  DFQD1 \mem_reg[207][9]  ( .D(n1350), .CP(clk), .Q(\mem[207][9] ) );
  DFQD1 \mem_reg[207][8]  ( .D(n1349), .CP(clk), .Q(\mem[207][8] ) );
  DFQD1 \mem_reg[207][7]  ( .D(n1348), .CP(clk), .Q(\mem[207][7] ) );
  DFQD1 \mem_reg[207][6]  ( .D(n1347), .CP(clk), .Q(\mem[207][6] ) );
  DFQD1 \mem_reg[207][5]  ( .D(n1346), .CP(clk), .Q(\mem[207][5] ) );
  DFQD1 \mem_reg[207][4]  ( .D(n1345), .CP(clk), .Q(\mem[207][4] ) );
  DFQD1 \mem_reg[207][3]  ( .D(n1344), .CP(clk), .Q(\mem[207][3] ) );
  DFQD1 \mem_reg[207][2]  ( .D(n1343), .CP(clk), .Q(\mem[207][2] ) );
  DFQD1 \mem_reg[207][1]  ( .D(n1342), .CP(clk), .Q(\mem[207][1] ) );
  DFQD1 \mem_reg[207][0]  ( .D(n1341), .CP(clk), .Q(\mem[207][0] ) );
  DFQD1 \mem_reg[208][15]  ( .D(n1340), .CP(clk), .Q(\mem[208][15] ) );
  DFQD1 \mem_reg[208][14]  ( .D(n1339), .CP(clk), .Q(\mem[208][14] ) );
  DFQD1 \mem_reg[208][13]  ( .D(n1338), .CP(clk), .Q(\mem[208][13] ) );
  DFQD1 \mem_reg[208][12]  ( .D(n1337), .CP(clk), .Q(\mem[208][12] ) );
  DFQD1 \mem_reg[208][11]  ( .D(n1336), .CP(clk), .Q(\mem[208][11] ) );
  DFQD1 \mem_reg[208][10]  ( .D(n1335), .CP(clk), .Q(\mem[208][10] ) );
  DFQD1 \mem_reg[208][9]  ( .D(n1334), .CP(clk), .Q(\mem[208][9] ) );
  DFQD1 \mem_reg[208][8]  ( .D(n1333), .CP(clk), .Q(\mem[208][8] ) );
  DFQD1 \mem_reg[208][7]  ( .D(n1332), .CP(clk), .Q(\mem[208][7] ) );
  DFQD1 \mem_reg[208][6]  ( .D(n1331), .CP(clk), .Q(\mem[208][6] ) );
  DFQD1 \mem_reg[208][5]  ( .D(n1330), .CP(clk), .Q(\mem[208][5] ) );
  DFQD1 \mem_reg[208][4]  ( .D(n1329), .CP(clk), .Q(\mem[208][4] ) );
  DFQD1 \mem_reg[208][3]  ( .D(n1328), .CP(clk), .Q(\mem[208][3] ) );
  DFQD1 \mem_reg[208][2]  ( .D(n1327), .CP(clk), .Q(\mem[208][2] ) );
  DFQD1 \mem_reg[208][1]  ( .D(n1326), .CP(clk), .Q(\mem[208][1] ) );
  DFQD1 \mem_reg[208][0]  ( .D(n1325), .CP(clk), .Q(\mem[208][0] ) );
  DFQD1 \mem_reg[209][15]  ( .D(n1324), .CP(clk), .Q(\mem[209][15] ) );
  DFQD1 \mem_reg[209][14]  ( .D(n1323), .CP(clk), .Q(\mem[209][14] ) );
  DFQD1 \mem_reg[209][13]  ( .D(n1322), .CP(clk), .Q(\mem[209][13] ) );
  DFQD1 \mem_reg[209][12]  ( .D(n1321), .CP(clk), .Q(\mem[209][12] ) );
  DFQD1 \mem_reg[209][11]  ( .D(n1320), .CP(clk), .Q(\mem[209][11] ) );
  DFQD1 \mem_reg[209][10]  ( .D(n1319), .CP(clk), .Q(\mem[209][10] ) );
  DFQD1 \mem_reg[209][9]  ( .D(n1318), .CP(clk), .Q(\mem[209][9] ) );
  DFQD1 \mem_reg[209][8]  ( .D(n1317), .CP(clk), .Q(\mem[209][8] ) );
  DFQD1 \mem_reg[209][7]  ( .D(n1316), .CP(clk), .Q(\mem[209][7] ) );
  DFQD1 \mem_reg[209][6]  ( .D(n1315), .CP(clk), .Q(\mem[209][6] ) );
  DFQD1 \mem_reg[209][5]  ( .D(n1314), .CP(clk), .Q(\mem[209][5] ) );
  DFQD1 \mem_reg[209][4]  ( .D(n1313), .CP(clk), .Q(\mem[209][4] ) );
  DFQD1 \mem_reg[209][3]  ( .D(n1312), .CP(clk), .Q(\mem[209][3] ) );
  DFQD1 \mem_reg[209][2]  ( .D(n1311), .CP(clk), .Q(\mem[209][2] ) );
  DFQD1 \mem_reg[209][1]  ( .D(n1310), .CP(clk), .Q(\mem[209][1] ) );
  DFQD1 \mem_reg[209][0]  ( .D(n1309), .CP(clk), .Q(\mem[209][0] ) );
  DFQD1 \mem_reg[210][15]  ( .D(n1308), .CP(clk), .Q(\mem[210][15] ) );
  DFQD1 \mem_reg[210][14]  ( .D(n1307), .CP(clk), .Q(\mem[210][14] ) );
  DFQD1 \mem_reg[210][13]  ( .D(n1306), .CP(clk), .Q(\mem[210][13] ) );
  DFQD1 \mem_reg[210][12]  ( .D(n1305), .CP(clk), .Q(\mem[210][12] ) );
  DFQD1 \mem_reg[210][11]  ( .D(n1304), .CP(clk), .Q(\mem[210][11] ) );
  DFQD1 \mem_reg[210][10]  ( .D(n1303), .CP(clk), .Q(\mem[210][10] ) );
  DFQD1 \mem_reg[210][9]  ( .D(n1302), .CP(clk), .Q(\mem[210][9] ) );
  DFQD1 \mem_reg[210][8]  ( .D(n1301), .CP(clk), .Q(\mem[210][8] ) );
  DFQD1 \mem_reg[210][7]  ( .D(n1300), .CP(clk), .Q(\mem[210][7] ) );
  DFQD1 \mem_reg[210][6]  ( .D(n1299), .CP(clk), .Q(\mem[210][6] ) );
  DFQD1 \mem_reg[210][5]  ( .D(n1298), .CP(clk), .Q(\mem[210][5] ) );
  DFQD1 \mem_reg[210][4]  ( .D(n1297), .CP(clk), .Q(\mem[210][4] ) );
  DFQD1 \mem_reg[210][3]  ( .D(n1296), .CP(clk), .Q(\mem[210][3] ) );
  DFQD1 \mem_reg[210][2]  ( .D(n1295), .CP(clk), .Q(\mem[210][2] ) );
  DFQD1 \mem_reg[210][1]  ( .D(n1294), .CP(clk), .Q(\mem[210][1] ) );
  DFQD1 \mem_reg[210][0]  ( .D(n1293), .CP(clk), .Q(\mem[210][0] ) );
  DFQD1 \mem_reg[211][15]  ( .D(n1292), .CP(clk), .Q(\mem[211][15] ) );
  DFQD1 \mem_reg[211][14]  ( .D(n1291), .CP(clk), .Q(\mem[211][14] ) );
  DFQD1 \mem_reg[211][13]  ( .D(n1290), .CP(clk), .Q(\mem[211][13] ) );
  DFQD1 \mem_reg[211][12]  ( .D(n1289), .CP(clk), .Q(\mem[211][12] ) );
  DFQD1 \mem_reg[211][11]  ( .D(n1288), .CP(clk), .Q(\mem[211][11] ) );
  DFQD1 \mem_reg[211][10]  ( .D(n1287), .CP(clk), .Q(\mem[211][10] ) );
  DFQD1 \mem_reg[211][9]  ( .D(n1286), .CP(clk), .Q(\mem[211][9] ) );
  DFQD1 \mem_reg[211][8]  ( .D(n1285), .CP(clk), .Q(\mem[211][8] ) );
  DFQD1 \mem_reg[211][7]  ( .D(n1284), .CP(clk), .Q(\mem[211][7] ) );
  DFQD1 \mem_reg[211][6]  ( .D(n1283), .CP(clk), .Q(\mem[211][6] ) );
  DFQD1 \mem_reg[211][5]  ( .D(n1282), .CP(clk), .Q(\mem[211][5] ) );
  DFQD1 \mem_reg[211][4]  ( .D(n1281), .CP(clk), .Q(\mem[211][4] ) );
  DFQD1 \mem_reg[211][3]  ( .D(n1280), .CP(clk), .Q(\mem[211][3] ) );
  DFQD1 \mem_reg[211][2]  ( .D(n1279), .CP(clk), .Q(\mem[211][2] ) );
  DFQD1 \mem_reg[211][1]  ( .D(n1278), .CP(clk), .Q(\mem[211][1] ) );
  DFQD1 \mem_reg[211][0]  ( .D(n1277), .CP(clk), .Q(\mem[211][0] ) );
  DFQD1 \mem_reg[212][15]  ( .D(n1276), .CP(clk), .Q(\mem[212][15] ) );
  DFQD1 \mem_reg[212][14]  ( .D(n1275), .CP(clk), .Q(\mem[212][14] ) );
  DFQD1 \mem_reg[212][13]  ( .D(n1274), .CP(clk), .Q(\mem[212][13] ) );
  DFQD1 \mem_reg[212][12]  ( .D(n1273), .CP(clk), .Q(\mem[212][12] ) );
  DFQD1 \mem_reg[212][11]  ( .D(n1272), .CP(clk), .Q(\mem[212][11] ) );
  DFQD1 \mem_reg[212][10]  ( .D(n1271), .CP(clk), .Q(\mem[212][10] ) );
  DFQD1 \mem_reg[212][9]  ( .D(n1270), .CP(clk), .Q(\mem[212][9] ) );
  DFQD1 \mem_reg[212][8]  ( .D(n1269), .CP(clk), .Q(\mem[212][8] ) );
  DFQD1 \mem_reg[212][7]  ( .D(n1268), .CP(clk), .Q(\mem[212][7] ) );
  DFQD1 \mem_reg[212][6]  ( .D(n1267), .CP(clk), .Q(\mem[212][6] ) );
  DFQD1 \mem_reg[212][5]  ( .D(n1266), .CP(clk), .Q(\mem[212][5] ) );
  DFQD1 \mem_reg[212][4]  ( .D(n1265), .CP(clk), .Q(\mem[212][4] ) );
  DFQD1 \mem_reg[212][3]  ( .D(n1264), .CP(clk), .Q(\mem[212][3] ) );
  DFQD1 \mem_reg[212][2]  ( .D(n1263), .CP(clk), .Q(\mem[212][2] ) );
  DFQD1 \mem_reg[212][1]  ( .D(n1262), .CP(clk), .Q(\mem[212][1] ) );
  DFQD1 \mem_reg[212][0]  ( .D(n1261), .CP(clk), .Q(\mem[212][0] ) );
  DFQD1 \mem_reg[213][15]  ( .D(n1260), .CP(clk), .Q(\mem[213][15] ) );
  DFQD1 \mem_reg[213][14]  ( .D(n1259), .CP(clk), .Q(\mem[213][14] ) );
  DFQD1 \mem_reg[213][13]  ( .D(n1258), .CP(clk), .Q(\mem[213][13] ) );
  DFQD1 \mem_reg[213][12]  ( .D(n1257), .CP(clk), .Q(\mem[213][12] ) );
  DFQD1 \mem_reg[213][11]  ( .D(n1256), .CP(clk), .Q(\mem[213][11] ) );
  DFQD1 \mem_reg[213][10]  ( .D(n1255), .CP(clk), .Q(\mem[213][10] ) );
  DFQD1 \mem_reg[213][9]  ( .D(n1254), .CP(clk), .Q(\mem[213][9] ) );
  DFQD1 \mem_reg[213][8]  ( .D(n1253), .CP(clk), .Q(\mem[213][8] ) );
  DFQD1 \mem_reg[213][7]  ( .D(n1252), .CP(clk), .Q(\mem[213][7] ) );
  DFQD1 \mem_reg[213][6]  ( .D(n1251), .CP(clk), .Q(\mem[213][6] ) );
  DFQD1 \mem_reg[213][5]  ( .D(n1250), .CP(clk), .Q(\mem[213][5] ) );
  DFQD1 \mem_reg[213][4]  ( .D(n1249), .CP(clk), .Q(\mem[213][4] ) );
  DFQD1 \mem_reg[213][3]  ( .D(n1248), .CP(clk), .Q(\mem[213][3] ) );
  DFQD1 \mem_reg[213][2]  ( .D(n1247), .CP(clk), .Q(\mem[213][2] ) );
  DFQD1 \mem_reg[213][1]  ( .D(n1246), .CP(clk), .Q(\mem[213][1] ) );
  DFQD1 \mem_reg[213][0]  ( .D(n1245), .CP(clk), .Q(\mem[213][0] ) );
  DFQD1 \mem_reg[214][15]  ( .D(n1244), .CP(clk), .Q(\mem[214][15] ) );
  DFQD1 \mem_reg[214][14]  ( .D(n1243), .CP(clk), .Q(\mem[214][14] ) );
  DFQD1 \mem_reg[214][13]  ( .D(n1242), .CP(clk), .Q(\mem[214][13] ) );
  DFQD1 \mem_reg[214][12]  ( .D(n1241), .CP(clk), .Q(\mem[214][12] ) );
  DFQD1 \mem_reg[214][11]  ( .D(n1240), .CP(clk), .Q(\mem[214][11] ) );
  DFQD1 \mem_reg[214][10]  ( .D(n1239), .CP(clk), .Q(\mem[214][10] ) );
  DFQD1 \mem_reg[214][9]  ( .D(n1238), .CP(clk), .Q(\mem[214][9] ) );
  DFQD1 \mem_reg[214][8]  ( .D(n1237), .CP(clk), .Q(\mem[214][8] ) );
  DFQD1 \mem_reg[214][7]  ( .D(n1236), .CP(clk), .Q(\mem[214][7] ) );
  DFQD1 \mem_reg[214][6]  ( .D(n1235), .CP(clk), .Q(\mem[214][6] ) );
  DFQD1 \mem_reg[214][5]  ( .D(n1234), .CP(clk), .Q(\mem[214][5] ) );
  DFQD1 \mem_reg[214][4]  ( .D(n1233), .CP(clk), .Q(\mem[214][4] ) );
  DFQD1 \mem_reg[214][3]  ( .D(n1232), .CP(clk), .Q(\mem[214][3] ) );
  DFQD1 \mem_reg[214][2]  ( .D(n1231), .CP(clk), .Q(\mem[214][2] ) );
  DFQD1 \mem_reg[214][1]  ( .D(n1230), .CP(clk), .Q(\mem[214][1] ) );
  DFQD1 \mem_reg[214][0]  ( .D(n1229), .CP(clk), .Q(\mem[214][0] ) );
  DFQD1 \mem_reg[215][15]  ( .D(n1228), .CP(clk), .Q(\mem[215][15] ) );
  DFQD1 \mem_reg[215][14]  ( .D(n1227), .CP(clk), .Q(\mem[215][14] ) );
  DFQD1 \mem_reg[215][13]  ( .D(n1226), .CP(clk), .Q(\mem[215][13] ) );
  DFQD1 \mem_reg[215][12]  ( .D(n1225), .CP(clk), .Q(\mem[215][12] ) );
  DFQD1 \mem_reg[215][11]  ( .D(n1224), .CP(clk), .Q(\mem[215][11] ) );
  DFQD1 \mem_reg[215][10]  ( .D(n1223), .CP(clk), .Q(\mem[215][10] ) );
  DFQD1 \mem_reg[215][9]  ( .D(n1222), .CP(clk), .Q(\mem[215][9] ) );
  DFQD1 \mem_reg[215][8]  ( .D(n1221), .CP(clk), .Q(\mem[215][8] ) );
  DFQD1 \mem_reg[215][7]  ( .D(n1220), .CP(clk), .Q(\mem[215][7] ) );
  DFQD1 \mem_reg[215][6]  ( .D(n1219), .CP(clk), .Q(\mem[215][6] ) );
  DFQD1 \mem_reg[215][5]  ( .D(n1218), .CP(clk), .Q(\mem[215][5] ) );
  DFQD1 \mem_reg[215][4]  ( .D(n1217), .CP(clk), .Q(\mem[215][4] ) );
  DFQD1 \mem_reg[215][3]  ( .D(n1216), .CP(clk), .Q(\mem[215][3] ) );
  DFQD1 \mem_reg[215][2]  ( .D(n1215), .CP(clk), .Q(\mem[215][2] ) );
  DFQD1 \mem_reg[215][1]  ( .D(n1214), .CP(clk), .Q(\mem[215][1] ) );
  DFQD1 \mem_reg[215][0]  ( .D(n1213), .CP(clk), .Q(\mem[215][0] ) );
  DFQD1 \mem_reg[216][15]  ( .D(n1212), .CP(clk), .Q(\mem[216][15] ) );
  DFQD1 \mem_reg[216][14]  ( .D(n1211), .CP(clk), .Q(\mem[216][14] ) );
  DFQD1 \mem_reg[216][13]  ( .D(n1210), .CP(clk), .Q(\mem[216][13] ) );
  DFQD1 \mem_reg[216][12]  ( .D(n1209), .CP(clk), .Q(\mem[216][12] ) );
  DFQD1 \mem_reg[216][11]  ( .D(n1208), .CP(clk), .Q(\mem[216][11] ) );
  DFQD1 \mem_reg[216][10]  ( .D(n1207), .CP(clk), .Q(\mem[216][10] ) );
  DFQD1 \mem_reg[216][9]  ( .D(n1206), .CP(clk), .Q(\mem[216][9] ) );
  DFQD1 \mem_reg[216][8]  ( .D(n1205), .CP(clk), .Q(\mem[216][8] ) );
  DFQD1 \mem_reg[216][7]  ( .D(n1204), .CP(clk), .Q(\mem[216][7] ) );
  DFQD1 \mem_reg[216][6]  ( .D(n1203), .CP(clk), .Q(\mem[216][6] ) );
  DFQD1 \mem_reg[216][5]  ( .D(n1202), .CP(clk), .Q(\mem[216][5] ) );
  DFQD1 \mem_reg[216][4]  ( .D(n1201), .CP(clk), .Q(\mem[216][4] ) );
  DFQD1 \mem_reg[216][3]  ( .D(n1200), .CP(clk), .Q(\mem[216][3] ) );
  DFQD1 \mem_reg[216][2]  ( .D(n1199), .CP(clk), .Q(\mem[216][2] ) );
  DFQD1 \mem_reg[216][1]  ( .D(n1198), .CP(clk), .Q(\mem[216][1] ) );
  DFQD1 \mem_reg[216][0]  ( .D(n1197), .CP(clk), .Q(\mem[216][0] ) );
  DFQD1 \mem_reg[217][15]  ( .D(n1196), .CP(clk), .Q(\mem[217][15] ) );
  DFQD1 \mem_reg[217][14]  ( .D(n1195), .CP(clk), .Q(\mem[217][14] ) );
  DFQD1 \mem_reg[217][13]  ( .D(n1194), .CP(clk), .Q(\mem[217][13] ) );
  DFQD1 \mem_reg[217][12]  ( .D(n1193), .CP(clk), .Q(\mem[217][12] ) );
  DFQD1 \mem_reg[217][11]  ( .D(n1192), .CP(clk), .Q(\mem[217][11] ) );
  DFQD1 \mem_reg[217][10]  ( .D(n1191), .CP(clk), .Q(\mem[217][10] ) );
  DFQD1 \mem_reg[217][9]  ( .D(n1190), .CP(clk), .Q(\mem[217][9] ) );
  DFQD1 \mem_reg[217][8]  ( .D(n1189), .CP(clk), .Q(\mem[217][8] ) );
  DFQD1 \mem_reg[217][7]  ( .D(n1188), .CP(clk), .Q(\mem[217][7] ) );
  DFQD1 \mem_reg[217][6]  ( .D(n1187), .CP(clk), .Q(\mem[217][6] ) );
  DFQD1 \mem_reg[217][5]  ( .D(n1186), .CP(clk), .Q(\mem[217][5] ) );
  DFQD1 \mem_reg[217][4]  ( .D(n1185), .CP(clk), .Q(\mem[217][4] ) );
  DFQD1 \mem_reg[217][3]  ( .D(n1184), .CP(clk), .Q(\mem[217][3] ) );
  DFQD1 \mem_reg[217][2]  ( .D(n1183), .CP(clk), .Q(\mem[217][2] ) );
  DFQD1 \mem_reg[217][1]  ( .D(n1182), .CP(clk), .Q(\mem[217][1] ) );
  DFQD1 \mem_reg[217][0]  ( .D(n1181), .CP(clk), .Q(\mem[217][0] ) );
  DFQD1 \mem_reg[218][15]  ( .D(n1180), .CP(clk), .Q(\mem[218][15] ) );
  DFQD1 \mem_reg[218][14]  ( .D(n1179), .CP(clk), .Q(\mem[218][14] ) );
  DFQD1 \mem_reg[218][13]  ( .D(n1178), .CP(clk), .Q(\mem[218][13] ) );
  DFQD1 \mem_reg[218][12]  ( .D(n1177), .CP(clk), .Q(\mem[218][12] ) );
  DFQD1 \mem_reg[218][11]  ( .D(n1176), .CP(clk), .Q(\mem[218][11] ) );
  DFQD1 \mem_reg[218][10]  ( .D(n1175), .CP(clk), .Q(\mem[218][10] ) );
  DFQD1 \mem_reg[218][9]  ( .D(n1174), .CP(clk), .Q(\mem[218][9] ) );
  DFQD1 \mem_reg[218][8]  ( .D(n1173), .CP(clk), .Q(\mem[218][8] ) );
  DFQD1 \mem_reg[218][7]  ( .D(n1172), .CP(clk), .Q(\mem[218][7] ) );
  DFQD1 \mem_reg[218][6]  ( .D(n1171), .CP(clk), .Q(\mem[218][6] ) );
  DFQD1 \mem_reg[218][5]  ( .D(n1170), .CP(clk), .Q(\mem[218][5] ) );
  DFQD1 \mem_reg[218][4]  ( .D(n1169), .CP(clk), .Q(\mem[218][4] ) );
  DFQD1 \mem_reg[218][3]  ( .D(n1168), .CP(clk), .Q(\mem[218][3] ) );
  DFQD1 \mem_reg[218][2]  ( .D(n1167), .CP(clk), .Q(\mem[218][2] ) );
  DFQD1 \mem_reg[218][1]  ( .D(n1166), .CP(clk), .Q(\mem[218][1] ) );
  DFQD1 \mem_reg[218][0]  ( .D(n1165), .CP(clk), .Q(\mem[218][0] ) );
  DFQD1 \mem_reg[219][15]  ( .D(n1164), .CP(clk), .Q(\mem[219][15] ) );
  DFQD1 \mem_reg[219][14]  ( .D(n1163), .CP(clk), .Q(\mem[219][14] ) );
  DFQD1 \mem_reg[219][13]  ( .D(n1162), .CP(clk), .Q(\mem[219][13] ) );
  DFQD1 \mem_reg[219][12]  ( .D(n1161), .CP(clk), .Q(\mem[219][12] ) );
  DFQD1 \mem_reg[219][11]  ( .D(n1160), .CP(clk), .Q(\mem[219][11] ) );
  DFQD1 \mem_reg[219][10]  ( .D(n1159), .CP(clk), .Q(\mem[219][10] ) );
  DFQD1 \mem_reg[219][9]  ( .D(n1158), .CP(clk), .Q(\mem[219][9] ) );
  DFQD1 \mem_reg[219][8]  ( .D(n1157), .CP(clk), .Q(\mem[219][8] ) );
  DFQD1 \mem_reg[219][7]  ( .D(n1156), .CP(clk), .Q(\mem[219][7] ) );
  DFQD1 \mem_reg[219][6]  ( .D(n1155), .CP(clk), .Q(\mem[219][6] ) );
  DFQD1 \mem_reg[219][5]  ( .D(n1154), .CP(clk), .Q(\mem[219][5] ) );
  DFQD1 \mem_reg[219][4]  ( .D(n1153), .CP(clk), .Q(\mem[219][4] ) );
  DFQD1 \mem_reg[219][3]  ( .D(n1152), .CP(clk), .Q(\mem[219][3] ) );
  DFQD1 \mem_reg[219][2]  ( .D(n1151), .CP(clk), .Q(\mem[219][2] ) );
  DFQD1 \mem_reg[219][1]  ( .D(n1150), .CP(clk), .Q(\mem[219][1] ) );
  DFQD1 \mem_reg[219][0]  ( .D(n1149), .CP(clk), .Q(\mem[219][0] ) );
  DFQD1 \mem_reg[220][15]  ( .D(n1148), .CP(clk), .Q(\mem[220][15] ) );
  DFQD1 \mem_reg[220][14]  ( .D(n1147), .CP(clk), .Q(\mem[220][14] ) );
  DFQD1 \mem_reg[220][13]  ( .D(n1146), .CP(clk), .Q(\mem[220][13] ) );
  DFQD1 \mem_reg[220][12]  ( .D(n1145), .CP(clk), .Q(\mem[220][12] ) );
  DFQD1 \mem_reg[220][11]  ( .D(n1144), .CP(clk), .Q(\mem[220][11] ) );
  DFQD1 \mem_reg[220][10]  ( .D(n1143), .CP(clk), .Q(\mem[220][10] ) );
  DFQD1 \mem_reg[220][9]  ( .D(n1142), .CP(clk), .Q(\mem[220][9] ) );
  DFQD1 \mem_reg[220][8]  ( .D(n1141), .CP(clk), .Q(\mem[220][8] ) );
  DFQD1 \mem_reg[220][7]  ( .D(n1140), .CP(clk), .Q(\mem[220][7] ) );
  DFQD1 \mem_reg[220][6]  ( .D(n1139), .CP(clk), .Q(\mem[220][6] ) );
  DFQD1 \mem_reg[220][5]  ( .D(n1138), .CP(clk), .Q(\mem[220][5] ) );
  DFQD1 \mem_reg[220][4]  ( .D(n1137), .CP(clk), .Q(\mem[220][4] ) );
  DFQD1 \mem_reg[220][3]  ( .D(n1136), .CP(clk), .Q(\mem[220][3] ) );
  DFQD1 \mem_reg[220][2]  ( .D(n1135), .CP(clk), .Q(\mem[220][2] ) );
  DFQD1 \mem_reg[220][1]  ( .D(n1134), .CP(clk), .Q(\mem[220][1] ) );
  DFQD1 \mem_reg[220][0]  ( .D(n1133), .CP(clk), .Q(\mem[220][0] ) );
  DFQD1 \mem_reg[221][15]  ( .D(n1132), .CP(clk), .Q(\mem[221][15] ) );
  DFQD1 \mem_reg[221][14]  ( .D(n1131), .CP(clk), .Q(\mem[221][14] ) );
  DFQD1 \mem_reg[221][13]  ( .D(n1130), .CP(clk), .Q(\mem[221][13] ) );
  DFQD1 \mem_reg[221][12]  ( .D(n1129), .CP(clk), .Q(\mem[221][12] ) );
  DFQD1 \mem_reg[221][11]  ( .D(n1128), .CP(clk), .Q(\mem[221][11] ) );
  DFQD1 \mem_reg[221][10]  ( .D(n1127), .CP(clk), .Q(\mem[221][10] ) );
  DFQD1 \mem_reg[221][9]  ( .D(n1126), .CP(clk), .Q(\mem[221][9] ) );
  DFQD1 \mem_reg[221][8]  ( .D(n1125), .CP(clk), .Q(\mem[221][8] ) );
  DFQD1 \mem_reg[221][7]  ( .D(n1124), .CP(clk), .Q(\mem[221][7] ) );
  DFQD1 \mem_reg[221][6]  ( .D(n1123), .CP(clk), .Q(\mem[221][6] ) );
  DFQD1 \mem_reg[221][5]  ( .D(n1122), .CP(clk), .Q(\mem[221][5] ) );
  DFQD1 \mem_reg[221][4]  ( .D(n1121), .CP(clk), .Q(\mem[221][4] ) );
  DFQD1 \mem_reg[221][3]  ( .D(n1120), .CP(clk), .Q(\mem[221][3] ) );
  DFQD1 \mem_reg[221][2]  ( .D(n1119), .CP(clk), .Q(\mem[221][2] ) );
  DFQD1 \mem_reg[221][1]  ( .D(n1118), .CP(clk), .Q(\mem[221][1] ) );
  DFQD1 \mem_reg[221][0]  ( .D(n1117), .CP(clk), .Q(\mem[221][0] ) );
  DFQD1 \mem_reg[222][15]  ( .D(n1116), .CP(clk), .Q(\mem[222][15] ) );
  DFQD1 \mem_reg[222][14]  ( .D(n1115), .CP(clk), .Q(\mem[222][14] ) );
  DFQD1 \mem_reg[222][13]  ( .D(n1114), .CP(clk), .Q(\mem[222][13] ) );
  DFQD1 \mem_reg[222][12]  ( .D(n1113), .CP(clk), .Q(\mem[222][12] ) );
  DFQD1 \mem_reg[222][11]  ( .D(n1112), .CP(clk), .Q(\mem[222][11] ) );
  DFQD1 \mem_reg[222][10]  ( .D(n1111), .CP(clk), .Q(\mem[222][10] ) );
  DFQD1 \mem_reg[222][9]  ( .D(n1110), .CP(clk), .Q(\mem[222][9] ) );
  DFQD1 \mem_reg[222][8]  ( .D(n1109), .CP(clk), .Q(\mem[222][8] ) );
  DFQD1 \mem_reg[222][7]  ( .D(n1108), .CP(clk), .Q(\mem[222][7] ) );
  DFQD1 \mem_reg[222][6]  ( .D(n1107), .CP(clk), .Q(\mem[222][6] ) );
  DFQD1 \mem_reg[222][5]  ( .D(n1106), .CP(clk), .Q(\mem[222][5] ) );
  DFQD1 \mem_reg[222][4]  ( .D(n1105), .CP(clk), .Q(\mem[222][4] ) );
  DFQD1 \mem_reg[222][3]  ( .D(n1104), .CP(clk), .Q(\mem[222][3] ) );
  DFQD1 \mem_reg[222][2]  ( .D(n1103), .CP(clk), .Q(\mem[222][2] ) );
  DFQD1 \mem_reg[222][1]  ( .D(n1102), .CP(clk), .Q(\mem[222][1] ) );
  DFQD1 \mem_reg[222][0]  ( .D(n1101), .CP(clk), .Q(\mem[222][0] ) );
  DFQD1 \mem_reg[223][15]  ( .D(n1100), .CP(clk), .Q(\mem[223][15] ) );
  DFQD1 \mem_reg[223][14]  ( .D(n1099), .CP(clk), .Q(\mem[223][14] ) );
  DFQD1 \mem_reg[223][13]  ( .D(n1098), .CP(clk), .Q(\mem[223][13] ) );
  DFQD1 \mem_reg[223][12]  ( .D(n1097), .CP(clk), .Q(\mem[223][12] ) );
  DFQD1 \mem_reg[223][11]  ( .D(n1096), .CP(clk), .Q(\mem[223][11] ) );
  DFQD1 \mem_reg[223][10]  ( .D(n1095), .CP(clk), .Q(\mem[223][10] ) );
  DFQD1 \mem_reg[223][9]  ( .D(n1094), .CP(clk), .Q(\mem[223][9] ) );
  DFQD1 \mem_reg[223][8]  ( .D(n1093), .CP(clk), .Q(\mem[223][8] ) );
  DFQD1 \mem_reg[223][7]  ( .D(n1092), .CP(clk), .Q(\mem[223][7] ) );
  DFQD1 \mem_reg[223][6]  ( .D(n1091), .CP(clk), .Q(\mem[223][6] ) );
  DFQD1 \mem_reg[223][5]  ( .D(n1090), .CP(clk), .Q(\mem[223][5] ) );
  DFQD1 \mem_reg[223][4]  ( .D(n1089), .CP(clk), .Q(\mem[223][4] ) );
  DFQD1 \mem_reg[223][3]  ( .D(n1088), .CP(clk), .Q(\mem[223][3] ) );
  DFQD1 \mem_reg[223][2]  ( .D(n1087), .CP(clk), .Q(\mem[223][2] ) );
  DFQD1 \mem_reg[223][1]  ( .D(n1086), .CP(clk), .Q(\mem[223][1] ) );
  DFQD1 \mem_reg[223][0]  ( .D(n1085), .CP(clk), .Q(\mem[223][0] ) );
  DFQD1 \mem_reg[224][15]  ( .D(n1084), .CP(clk), .Q(\mem[224][15] ) );
  DFQD1 \mem_reg[224][14]  ( .D(n1083), .CP(clk), .Q(\mem[224][14] ) );
  DFQD1 \mem_reg[224][13]  ( .D(n1082), .CP(clk), .Q(\mem[224][13] ) );
  DFQD1 \mem_reg[224][12]  ( .D(n1081), .CP(clk), .Q(\mem[224][12] ) );
  DFQD1 \mem_reg[224][11]  ( .D(n1080), .CP(clk), .Q(\mem[224][11] ) );
  DFQD1 \mem_reg[224][10]  ( .D(n1079), .CP(clk), .Q(\mem[224][10] ) );
  DFQD1 \mem_reg[224][9]  ( .D(n1078), .CP(clk), .Q(\mem[224][9] ) );
  DFQD1 \mem_reg[224][8]  ( .D(n1077), .CP(clk), .Q(\mem[224][8] ) );
  DFQD1 \mem_reg[224][7]  ( .D(n1076), .CP(clk), .Q(\mem[224][7] ) );
  DFQD1 \mem_reg[224][6]  ( .D(n1075), .CP(clk), .Q(\mem[224][6] ) );
  DFQD1 \mem_reg[224][5]  ( .D(n1074), .CP(clk), .Q(\mem[224][5] ) );
  DFQD1 \mem_reg[224][4]  ( .D(n1073), .CP(clk), .Q(\mem[224][4] ) );
  DFQD1 \mem_reg[224][3]  ( .D(n1072), .CP(clk), .Q(\mem[224][3] ) );
  DFQD1 \mem_reg[224][2]  ( .D(n1071), .CP(clk), .Q(\mem[224][2] ) );
  DFQD1 \mem_reg[224][1]  ( .D(n1070), .CP(clk), .Q(\mem[224][1] ) );
  DFQD1 \mem_reg[224][0]  ( .D(n1069), .CP(clk), .Q(\mem[224][0] ) );
  DFQD1 \mem_reg[225][15]  ( .D(n1068), .CP(clk), .Q(\mem[225][15] ) );
  DFQD1 \mem_reg[225][14]  ( .D(n1067), .CP(clk), .Q(\mem[225][14] ) );
  DFQD1 \mem_reg[225][13]  ( .D(n1066), .CP(clk), .Q(\mem[225][13] ) );
  DFQD1 \mem_reg[225][12]  ( .D(n1065), .CP(clk), .Q(\mem[225][12] ) );
  DFQD1 \mem_reg[225][11]  ( .D(n1064), .CP(clk), .Q(\mem[225][11] ) );
  DFQD1 \mem_reg[225][10]  ( .D(n1063), .CP(clk), .Q(\mem[225][10] ) );
  DFQD1 \mem_reg[225][9]  ( .D(n1062), .CP(clk), .Q(\mem[225][9] ) );
  DFQD1 \mem_reg[225][8]  ( .D(n1061), .CP(clk), .Q(\mem[225][8] ) );
  DFQD1 \mem_reg[225][7]  ( .D(n1060), .CP(clk), .Q(\mem[225][7] ) );
  DFQD1 \mem_reg[225][6]  ( .D(n1059), .CP(clk), .Q(\mem[225][6] ) );
  DFQD1 \mem_reg[225][5]  ( .D(n1058), .CP(clk), .Q(\mem[225][5] ) );
  DFQD1 \mem_reg[225][4]  ( .D(n1057), .CP(clk), .Q(\mem[225][4] ) );
  DFQD1 \mem_reg[225][3]  ( .D(n1056), .CP(clk), .Q(\mem[225][3] ) );
  DFQD1 \mem_reg[225][2]  ( .D(n1055), .CP(clk), .Q(\mem[225][2] ) );
  DFQD1 \mem_reg[225][1]  ( .D(n1054), .CP(clk), .Q(\mem[225][1] ) );
  DFQD1 \mem_reg[225][0]  ( .D(n1053), .CP(clk), .Q(\mem[225][0] ) );
  DFQD1 \mem_reg[226][15]  ( .D(n1052), .CP(clk), .Q(\mem[226][15] ) );
  DFQD1 \mem_reg[226][14]  ( .D(n1051), .CP(clk), .Q(\mem[226][14] ) );
  DFQD1 \mem_reg[226][13]  ( .D(n1050), .CP(clk), .Q(\mem[226][13] ) );
  DFQD1 \mem_reg[226][12]  ( .D(n1049), .CP(clk), .Q(\mem[226][12] ) );
  DFQD1 \mem_reg[226][11]  ( .D(n1048), .CP(clk), .Q(\mem[226][11] ) );
  DFQD1 \mem_reg[226][10]  ( .D(n1047), .CP(clk), .Q(\mem[226][10] ) );
  DFQD1 \mem_reg[226][9]  ( .D(n1046), .CP(clk), .Q(\mem[226][9] ) );
  DFQD1 \mem_reg[226][8]  ( .D(n1045), .CP(clk), .Q(\mem[226][8] ) );
  DFQD1 \mem_reg[226][7]  ( .D(n1044), .CP(clk), .Q(\mem[226][7] ) );
  DFQD1 \mem_reg[226][6]  ( .D(n1043), .CP(clk), .Q(\mem[226][6] ) );
  DFQD1 \mem_reg[226][5]  ( .D(n1042), .CP(clk), .Q(\mem[226][5] ) );
  DFQD1 \mem_reg[226][4]  ( .D(n1041), .CP(clk), .Q(\mem[226][4] ) );
  DFQD1 \mem_reg[226][3]  ( .D(n1040), .CP(clk), .Q(\mem[226][3] ) );
  DFQD1 \mem_reg[226][2]  ( .D(n1039), .CP(clk), .Q(\mem[226][2] ) );
  DFQD1 \mem_reg[226][1]  ( .D(n1038), .CP(clk), .Q(\mem[226][1] ) );
  DFQD1 \mem_reg[226][0]  ( .D(n1037), .CP(clk), .Q(\mem[226][0] ) );
  DFQD1 \mem_reg[227][15]  ( .D(n1036), .CP(clk), .Q(\mem[227][15] ) );
  DFQD1 \mem_reg[227][14]  ( .D(n1035), .CP(clk), .Q(\mem[227][14] ) );
  DFQD1 \mem_reg[227][13]  ( .D(n1034), .CP(clk), .Q(\mem[227][13] ) );
  DFQD1 \mem_reg[227][12]  ( .D(n1033), .CP(clk), .Q(\mem[227][12] ) );
  DFQD1 \mem_reg[227][11]  ( .D(n1032), .CP(clk), .Q(\mem[227][11] ) );
  DFQD1 \mem_reg[227][10]  ( .D(n1031), .CP(clk), .Q(\mem[227][10] ) );
  DFQD1 \mem_reg[227][9]  ( .D(n1030), .CP(clk), .Q(\mem[227][9] ) );
  DFQD1 \mem_reg[227][8]  ( .D(n1029), .CP(clk), .Q(\mem[227][8] ) );
  DFQD1 \mem_reg[227][7]  ( .D(n1028), .CP(clk), .Q(\mem[227][7] ) );
  DFQD1 \mem_reg[227][6]  ( .D(n1027), .CP(clk), .Q(\mem[227][6] ) );
  DFQD1 \mem_reg[227][5]  ( .D(n1026), .CP(clk), .Q(\mem[227][5] ) );
  DFQD1 \mem_reg[227][4]  ( .D(n1025), .CP(clk), .Q(\mem[227][4] ) );
  DFQD1 \mem_reg[227][3]  ( .D(n1024), .CP(clk), .Q(\mem[227][3] ) );
  DFQD1 \mem_reg[227][2]  ( .D(n1023), .CP(clk), .Q(\mem[227][2] ) );
  DFQD1 \mem_reg[227][1]  ( .D(n1022), .CP(clk), .Q(\mem[227][1] ) );
  DFQD1 \mem_reg[227][0]  ( .D(n1021), .CP(clk), .Q(\mem[227][0] ) );
  DFQD1 \mem_reg[228][15]  ( .D(n1020), .CP(clk), .Q(\mem[228][15] ) );
  DFQD1 \mem_reg[228][14]  ( .D(n1019), .CP(clk), .Q(\mem[228][14] ) );
  DFQD1 \mem_reg[228][13]  ( .D(n1018), .CP(clk), .Q(\mem[228][13] ) );
  DFQD1 \mem_reg[228][12]  ( .D(n1017), .CP(clk), .Q(\mem[228][12] ) );
  DFQD1 \mem_reg[228][11]  ( .D(n1016), .CP(clk), .Q(\mem[228][11] ) );
  DFQD1 \mem_reg[228][10]  ( .D(n1015), .CP(clk), .Q(\mem[228][10] ) );
  DFQD1 \mem_reg[228][9]  ( .D(n1014), .CP(clk), .Q(\mem[228][9] ) );
  DFQD1 \mem_reg[228][8]  ( .D(n1013), .CP(clk), .Q(\mem[228][8] ) );
  DFQD1 \mem_reg[228][7]  ( .D(n1012), .CP(clk), .Q(\mem[228][7] ) );
  DFQD1 \mem_reg[228][6]  ( .D(n1011), .CP(clk), .Q(\mem[228][6] ) );
  DFQD1 \mem_reg[228][5]  ( .D(n1010), .CP(clk), .Q(\mem[228][5] ) );
  DFQD1 \mem_reg[228][4]  ( .D(n1009), .CP(clk), .Q(\mem[228][4] ) );
  DFQD1 \mem_reg[228][3]  ( .D(n1008), .CP(clk), .Q(\mem[228][3] ) );
  DFQD1 \mem_reg[228][2]  ( .D(n1007), .CP(clk), .Q(\mem[228][2] ) );
  DFQD1 \mem_reg[228][1]  ( .D(n1006), .CP(clk), .Q(\mem[228][1] ) );
  DFQD1 \mem_reg[228][0]  ( .D(n1005), .CP(clk), .Q(\mem[228][0] ) );
  DFQD1 \mem_reg[229][15]  ( .D(n1004), .CP(clk), .Q(\mem[229][15] ) );
  DFQD1 \mem_reg[229][14]  ( .D(n1003), .CP(clk), .Q(\mem[229][14] ) );
  DFQD1 \mem_reg[229][13]  ( .D(n1002), .CP(clk), .Q(\mem[229][13] ) );
  DFQD1 \mem_reg[229][12]  ( .D(n1001), .CP(clk), .Q(\mem[229][12] ) );
  DFQD1 \mem_reg[229][11]  ( .D(n1000), .CP(clk), .Q(\mem[229][11] ) );
  DFQD1 \mem_reg[229][10]  ( .D(n999), .CP(clk), .Q(\mem[229][10] ) );
  DFQD1 \mem_reg[229][9]  ( .D(n998), .CP(clk), .Q(\mem[229][9] ) );
  DFQD1 \mem_reg[229][8]  ( .D(n997), .CP(clk), .Q(\mem[229][8] ) );
  DFQD1 \mem_reg[229][7]  ( .D(n996), .CP(clk), .Q(\mem[229][7] ) );
  DFQD1 \mem_reg[229][6]  ( .D(n995), .CP(clk), .Q(\mem[229][6] ) );
  DFQD1 \mem_reg[229][5]  ( .D(n994), .CP(clk), .Q(\mem[229][5] ) );
  DFQD1 \mem_reg[229][4]  ( .D(n993), .CP(clk), .Q(\mem[229][4] ) );
  DFQD1 \mem_reg[229][3]  ( .D(n992), .CP(clk), .Q(\mem[229][3] ) );
  DFQD1 \mem_reg[229][2]  ( .D(n991), .CP(clk), .Q(\mem[229][2] ) );
  DFQD1 \mem_reg[229][1]  ( .D(n990), .CP(clk), .Q(\mem[229][1] ) );
  DFQD1 \mem_reg[229][0]  ( .D(n989), .CP(clk), .Q(\mem[229][0] ) );
  DFQD1 \mem_reg[230][15]  ( .D(n988), .CP(clk), .Q(\mem[230][15] ) );
  DFQD1 \mem_reg[230][14]  ( .D(n987), .CP(clk), .Q(\mem[230][14] ) );
  DFQD1 \mem_reg[230][13]  ( .D(n986), .CP(clk), .Q(\mem[230][13] ) );
  DFQD1 \mem_reg[230][12]  ( .D(n985), .CP(clk), .Q(\mem[230][12] ) );
  DFQD1 \mem_reg[230][11]  ( .D(n984), .CP(clk), .Q(\mem[230][11] ) );
  DFQD1 \mem_reg[230][10]  ( .D(n983), .CP(clk), .Q(\mem[230][10] ) );
  DFQD1 \mem_reg[230][9]  ( .D(n982), .CP(clk), .Q(\mem[230][9] ) );
  DFQD1 \mem_reg[230][8]  ( .D(n981), .CP(clk), .Q(\mem[230][8] ) );
  DFQD1 \mem_reg[230][7]  ( .D(n980), .CP(clk), .Q(\mem[230][7] ) );
  DFQD1 \mem_reg[230][6]  ( .D(n979), .CP(clk), .Q(\mem[230][6] ) );
  DFQD1 \mem_reg[230][5]  ( .D(n978), .CP(clk), .Q(\mem[230][5] ) );
  DFQD1 \mem_reg[230][4]  ( .D(n977), .CP(clk), .Q(\mem[230][4] ) );
  DFQD1 \mem_reg[230][3]  ( .D(n976), .CP(clk), .Q(\mem[230][3] ) );
  DFQD1 \mem_reg[230][2]  ( .D(n975), .CP(clk), .Q(\mem[230][2] ) );
  DFQD1 \mem_reg[230][1]  ( .D(n974), .CP(clk), .Q(\mem[230][1] ) );
  DFQD1 \mem_reg[230][0]  ( .D(n973), .CP(clk), .Q(\mem[230][0] ) );
  DFQD1 \mem_reg[231][15]  ( .D(n972), .CP(clk), .Q(\mem[231][15] ) );
  DFQD1 \mem_reg[231][14]  ( .D(n971), .CP(clk), .Q(\mem[231][14] ) );
  DFQD1 \mem_reg[231][13]  ( .D(n970), .CP(clk), .Q(\mem[231][13] ) );
  DFQD1 \mem_reg[231][12]  ( .D(n969), .CP(clk), .Q(\mem[231][12] ) );
  DFQD1 \mem_reg[231][11]  ( .D(n968), .CP(clk), .Q(\mem[231][11] ) );
  DFQD1 \mem_reg[231][10]  ( .D(n967), .CP(clk), .Q(\mem[231][10] ) );
  DFQD1 \mem_reg[231][9]  ( .D(n966), .CP(clk), .Q(\mem[231][9] ) );
  DFQD1 \mem_reg[231][8]  ( .D(n965), .CP(clk), .Q(\mem[231][8] ) );
  DFQD1 \mem_reg[231][7]  ( .D(n964), .CP(clk), .Q(\mem[231][7] ) );
  DFQD1 \mem_reg[231][6]  ( .D(n963), .CP(clk), .Q(\mem[231][6] ) );
  DFQD1 \mem_reg[231][5]  ( .D(n962), .CP(clk), .Q(\mem[231][5] ) );
  DFQD1 \mem_reg[231][4]  ( .D(n961), .CP(clk), .Q(\mem[231][4] ) );
  DFQD1 \mem_reg[231][3]  ( .D(n960), .CP(clk), .Q(\mem[231][3] ) );
  DFQD1 \mem_reg[231][2]  ( .D(n959), .CP(clk), .Q(\mem[231][2] ) );
  DFQD1 \mem_reg[231][1]  ( .D(n958), .CP(clk), .Q(\mem[231][1] ) );
  DFQD1 \mem_reg[231][0]  ( .D(n957), .CP(clk), .Q(\mem[231][0] ) );
  DFQD1 \mem_reg[232][15]  ( .D(n956), .CP(clk), .Q(\mem[232][15] ) );
  DFQD1 \mem_reg[232][14]  ( .D(n955), .CP(clk), .Q(\mem[232][14] ) );
  DFQD1 \mem_reg[232][13]  ( .D(n954), .CP(clk), .Q(\mem[232][13] ) );
  DFQD1 \mem_reg[232][12]  ( .D(n953), .CP(clk), .Q(\mem[232][12] ) );
  DFQD1 \mem_reg[232][11]  ( .D(n952), .CP(clk), .Q(\mem[232][11] ) );
  DFQD1 \mem_reg[232][10]  ( .D(n951), .CP(clk), .Q(\mem[232][10] ) );
  DFQD1 \mem_reg[232][9]  ( .D(n950), .CP(clk), .Q(\mem[232][9] ) );
  DFQD1 \mem_reg[232][8]  ( .D(n949), .CP(clk), .Q(\mem[232][8] ) );
  DFQD1 \mem_reg[232][7]  ( .D(n948), .CP(clk), .Q(\mem[232][7] ) );
  DFQD1 \mem_reg[232][6]  ( .D(n947), .CP(clk), .Q(\mem[232][6] ) );
  DFQD1 \mem_reg[232][5]  ( .D(n946), .CP(clk), .Q(\mem[232][5] ) );
  DFQD1 \mem_reg[232][4]  ( .D(n945), .CP(clk), .Q(\mem[232][4] ) );
  DFQD1 \mem_reg[232][3]  ( .D(n944), .CP(clk), .Q(\mem[232][3] ) );
  DFQD1 \mem_reg[232][2]  ( .D(n943), .CP(clk), .Q(\mem[232][2] ) );
  DFQD1 \mem_reg[232][1]  ( .D(n942), .CP(clk), .Q(\mem[232][1] ) );
  DFQD1 \mem_reg[232][0]  ( .D(n941), .CP(clk), .Q(\mem[232][0] ) );
  DFQD1 \mem_reg[233][15]  ( .D(n940), .CP(clk), .Q(\mem[233][15] ) );
  DFQD1 \mem_reg[233][14]  ( .D(n939), .CP(clk), .Q(\mem[233][14] ) );
  DFQD1 \mem_reg[233][13]  ( .D(n938), .CP(clk), .Q(\mem[233][13] ) );
  DFQD1 \mem_reg[233][12]  ( .D(n937), .CP(clk), .Q(\mem[233][12] ) );
  DFQD1 \mem_reg[233][11]  ( .D(n936), .CP(clk), .Q(\mem[233][11] ) );
  DFQD1 \mem_reg[233][10]  ( .D(n935), .CP(clk), .Q(\mem[233][10] ) );
  DFQD1 \mem_reg[233][9]  ( .D(n934), .CP(clk), .Q(\mem[233][9] ) );
  DFQD1 \mem_reg[233][8]  ( .D(n933), .CP(clk), .Q(\mem[233][8] ) );
  DFQD1 \mem_reg[233][7]  ( .D(n932), .CP(clk), .Q(\mem[233][7] ) );
  DFQD1 \mem_reg[233][6]  ( .D(n931), .CP(clk), .Q(\mem[233][6] ) );
  DFQD1 \mem_reg[233][5]  ( .D(n930), .CP(clk), .Q(\mem[233][5] ) );
  DFQD1 \mem_reg[233][4]  ( .D(n929), .CP(clk), .Q(\mem[233][4] ) );
  DFQD1 \mem_reg[233][3]  ( .D(n928), .CP(clk), .Q(\mem[233][3] ) );
  DFQD1 \mem_reg[233][2]  ( .D(n927), .CP(clk), .Q(\mem[233][2] ) );
  DFQD1 \mem_reg[233][1]  ( .D(n926), .CP(clk), .Q(\mem[233][1] ) );
  DFQD1 \mem_reg[233][0]  ( .D(n925), .CP(clk), .Q(\mem[233][0] ) );
  DFQD1 \mem_reg[234][15]  ( .D(n924), .CP(clk), .Q(\mem[234][15] ) );
  DFQD1 \mem_reg[234][14]  ( .D(n923), .CP(clk), .Q(\mem[234][14] ) );
  DFQD1 \mem_reg[234][13]  ( .D(n922), .CP(clk), .Q(\mem[234][13] ) );
  DFQD1 \mem_reg[234][12]  ( .D(n921), .CP(clk), .Q(\mem[234][12] ) );
  DFQD1 \mem_reg[234][11]  ( .D(n920), .CP(clk), .Q(\mem[234][11] ) );
  DFQD1 \mem_reg[234][10]  ( .D(n919), .CP(clk), .Q(\mem[234][10] ) );
  DFQD1 \mem_reg[234][9]  ( .D(n918), .CP(clk), .Q(\mem[234][9] ) );
  DFQD1 \mem_reg[234][8]  ( .D(n917), .CP(clk), .Q(\mem[234][8] ) );
  DFQD1 \mem_reg[234][7]  ( .D(n916), .CP(clk), .Q(\mem[234][7] ) );
  DFQD1 \mem_reg[234][6]  ( .D(n915), .CP(clk), .Q(\mem[234][6] ) );
  DFQD1 \mem_reg[234][5]  ( .D(n914), .CP(clk), .Q(\mem[234][5] ) );
  DFQD1 \mem_reg[234][4]  ( .D(n913), .CP(clk), .Q(\mem[234][4] ) );
  DFQD1 \mem_reg[234][3]  ( .D(n912), .CP(clk), .Q(\mem[234][3] ) );
  DFQD1 \mem_reg[234][2]  ( .D(n911), .CP(clk), .Q(\mem[234][2] ) );
  DFQD1 \mem_reg[234][1]  ( .D(n910), .CP(clk), .Q(\mem[234][1] ) );
  DFQD1 \mem_reg[234][0]  ( .D(n909), .CP(clk), .Q(\mem[234][0] ) );
  DFQD1 \mem_reg[235][15]  ( .D(n908), .CP(clk), .Q(\mem[235][15] ) );
  DFQD1 \mem_reg[235][14]  ( .D(n907), .CP(clk), .Q(\mem[235][14] ) );
  DFQD1 \mem_reg[235][13]  ( .D(n906), .CP(clk), .Q(\mem[235][13] ) );
  DFQD1 \mem_reg[235][12]  ( .D(n905), .CP(clk), .Q(\mem[235][12] ) );
  DFQD1 \mem_reg[235][11]  ( .D(n904), .CP(clk), .Q(\mem[235][11] ) );
  DFQD1 \mem_reg[235][10]  ( .D(n903), .CP(clk), .Q(\mem[235][10] ) );
  DFQD1 \mem_reg[235][9]  ( .D(n902), .CP(clk), .Q(\mem[235][9] ) );
  DFQD1 \mem_reg[235][8]  ( .D(n901), .CP(clk), .Q(\mem[235][8] ) );
  DFQD1 \mem_reg[235][7]  ( .D(n900), .CP(clk), .Q(\mem[235][7] ) );
  DFQD1 \mem_reg[235][6]  ( .D(n899), .CP(clk), .Q(\mem[235][6] ) );
  DFQD1 \mem_reg[235][5]  ( .D(n898), .CP(clk), .Q(\mem[235][5] ) );
  DFQD1 \mem_reg[235][4]  ( .D(n897), .CP(clk), .Q(\mem[235][4] ) );
  DFQD1 \mem_reg[235][3]  ( .D(n896), .CP(clk), .Q(\mem[235][3] ) );
  DFQD1 \mem_reg[235][2]  ( .D(n895), .CP(clk), .Q(\mem[235][2] ) );
  DFQD1 \mem_reg[235][1]  ( .D(n894), .CP(clk), .Q(\mem[235][1] ) );
  DFQD1 \mem_reg[235][0]  ( .D(n893), .CP(clk), .Q(\mem[235][0] ) );
  DFQD1 \mem_reg[236][15]  ( .D(n892), .CP(clk), .Q(\mem[236][15] ) );
  DFQD1 \mem_reg[236][14]  ( .D(n891), .CP(clk), .Q(\mem[236][14] ) );
  DFQD1 \mem_reg[236][13]  ( .D(n890), .CP(clk), .Q(\mem[236][13] ) );
  DFQD1 \mem_reg[236][12]  ( .D(n889), .CP(clk), .Q(\mem[236][12] ) );
  DFQD1 \mem_reg[236][11]  ( .D(n888), .CP(clk), .Q(\mem[236][11] ) );
  DFQD1 \mem_reg[236][10]  ( .D(n887), .CP(clk), .Q(\mem[236][10] ) );
  DFQD1 \mem_reg[236][9]  ( .D(n886), .CP(clk), .Q(\mem[236][9] ) );
  DFQD1 \mem_reg[236][8]  ( .D(n885), .CP(clk), .Q(\mem[236][8] ) );
  DFQD1 \mem_reg[236][7]  ( .D(n884), .CP(clk), .Q(\mem[236][7] ) );
  DFQD1 \mem_reg[236][6]  ( .D(n883), .CP(clk), .Q(\mem[236][6] ) );
  DFQD1 \mem_reg[236][5]  ( .D(n882), .CP(clk), .Q(\mem[236][5] ) );
  DFQD1 \mem_reg[236][4]  ( .D(n881), .CP(clk), .Q(\mem[236][4] ) );
  DFQD1 \mem_reg[236][3]  ( .D(n880), .CP(clk), .Q(\mem[236][3] ) );
  DFQD1 \mem_reg[236][2]  ( .D(n879), .CP(clk), .Q(\mem[236][2] ) );
  DFQD1 \mem_reg[236][1]  ( .D(n878), .CP(clk), .Q(\mem[236][1] ) );
  DFQD1 \mem_reg[236][0]  ( .D(n877), .CP(clk), .Q(\mem[236][0] ) );
  DFQD1 \mem_reg[237][15]  ( .D(n876), .CP(clk), .Q(\mem[237][15] ) );
  DFQD1 \mem_reg[237][14]  ( .D(n875), .CP(clk), .Q(\mem[237][14] ) );
  DFQD1 \mem_reg[237][13]  ( .D(n874), .CP(clk), .Q(\mem[237][13] ) );
  DFQD1 \mem_reg[237][12]  ( .D(n873), .CP(clk), .Q(\mem[237][12] ) );
  DFQD1 \mem_reg[237][11]  ( .D(n872), .CP(clk), .Q(\mem[237][11] ) );
  DFQD1 \mem_reg[237][10]  ( .D(n871), .CP(clk), .Q(\mem[237][10] ) );
  DFQD1 \mem_reg[237][9]  ( .D(n870), .CP(clk), .Q(\mem[237][9] ) );
  DFQD1 \mem_reg[237][8]  ( .D(n869), .CP(clk), .Q(\mem[237][8] ) );
  DFQD1 \mem_reg[237][7]  ( .D(n868), .CP(clk), .Q(\mem[237][7] ) );
  DFQD1 \mem_reg[237][6]  ( .D(n867), .CP(clk), .Q(\mem[237][6] ) );
  DFQD1 \mem_reg[237][5]  ( .D(n866), .CP(clk), .Q(\mem[237][5] ) );
  DFQD1 \mem_reg[237][4]  ( .D(n865), .CP(clk), .Q(\mem[237][4] ) );
  DFQD1 \mem_reg[237][3]  ( .D(n864), .CP(clk), .Q(\mem[237][3] ) );
  DFQD1 \mem_reg[237][2]  ( .D(n863), .CP(clk), .Q(\mem[237][2] ) );
  DFQD1 \mem_reg[237][1]  ( .D(n862), .CP(clk), .Q(\mem[237][1] ) );
  DFQD1 \mem_reg[237][0]  ( .D(n861), .CP(clk), .Q(\mem[237][0] ) );
  DFQD1 \mem_reg[238][15]  ( .D(n860), .CP(clk), .Q(\mem[238][15] ) );
  DFQD1 \mem_reg[238][14]  ( .D(n859), .CP(clk), .Q(\mem[238][14] ) );
  DFQD1 \mem_reg[238][13]  ( .D(n858), .CP(clk), .Q(\mem[238][13] ) );
  DFQD1 \mem_reg[238][12]  ( .D(n857), .CP(clk), .Q(\mem[238][12] ) );
  DFQD1 \mem_reg[238][11]  ( .D(n856), .CP(clk), .Q(\mem[238][11] ) );
  DFQD1 \mem_reg[238][10]  ( .D(n855), .CP(clk), .Q(\mem[238][10] ) );
  DFQD1 \mem_reg[238][9]  ( .D(n854), .CP(clk), .Q(\mem[238][9] ) );
  DFQD1 \mem_reg[238][8]  ( .D(n853), .CP(clk), .Q(\mem[238][8] ) );
  DFQD1 \mem_reg[238][7]  ( .D(n852), .CP(clk), .Q(\mem[238][7] ) );
  DFQD1 \mem_reg[238][6]  ( .D(n851), .CP(clk), .Q(\mem[238][6] ) );
  DFQD1 \mem_reg[238][5]  ( .D(n850), .CP(clk), .Q(\mem[238][5] ) );
  DFQD1 \mem_reg[238][4]  ( .D(n849), .CP(clk), .Q(\mem[238][4] ) );
  DFQD1 \mem_reg[238][3]  ( .D(n848), .CP(clk), .Q(\mem[238][3] ) );
  DFQD1 \mem_reg[238][2]  ( .D(n847), .CP(clk), .Q(\mem[238][2] ) );
  DFQD1 \mem_reg[238][1]  ( .D(n846), .CP(clk), .Q(\mem[238][1] ) );
  DFQD1 \mem_reg[238][0]  ( .D(n845), .CP(clk), .Q(\mem[238][0] ) );
  DFQD1 \mem_reg[239][15]  ( .D(n844), .CP(clk), .Q(\mem[239][15] ) );
  DFQD1 \mem_reg[239][14]  ( .D(n843), .CP(clk), .Q(\mem[239][14] ) );
  DFQD1 \mem_reg[239][13]  ( .D(n842), .CP(clk), .Q(\mem[239][13] ) );
  DFQD1 \mem_reg[239][12]  ( .D(n841), .CP(clk), .Q(\mem[239][12] ) );
  DFQD1 \mem_reg[239][11]  ( .D(n840), .CP(clk), .Q(\mem[239][11] ) );
  DFQD1 \mem_reg[239][10]  ( .D(n839), .CP(clk), .Q(\mem[239][10] ) );
  DFQD1 \mem_reg[239][9]  ( .D(n838), .CP(clk), .Q(\mem[239][9] ) );
  DFQD1 \mem_reg[239][8]  ( .D(n837), .CP(clk), .Q(\mem[239][8] ) );
  DFQD1 \mem_reg[239][7]  ( .D(n836), .CP(clk), .Q(\mem[239][7] ) );
  DFQD1 \mem_reg[239][6]  ( .D(n835), .CP(clk), .Q(\mem[239][6] ) );
  DFQD1 \mem_reg[239][5]  ( .D(n834), .CP(clk), .Q(\mem[239][5] ) );
  DFQD1 \mem_reg[239][4]  ( .D(n833), .CP(clk), .Q(\mem[239][4] ) );
  DFQD1 \mem_reg[239][3]  ( .D(n832), .CP(clk), .Q(\mem[239][3] ) );
  DFQD1 \mem_reg[239][2]  ( .D(n831), .CP(clk), .Q(\mem[239][2] ) );
  DFQD1 \mem_reg[239][1]  ( .D(n830), .CP(clk), .Q(\mem[239][1] ) );
  DFQD1 \mem_reg[239][0]  ( .D(n829), .CP(clk), .Q(\mem[239][0] ) );
  DFQD1 \mem_reg[240][15]  ( .D(n828), .CP(clk), .Q(\mem[240][15] ) );
  DFQD1 \mem_reg[240][14]  ( .D(n827), .CP(clk), .Q(\mem[240][14] ) );
  DFQD1 \mem_reg[240][13]  ( .D(n826), .CP(clk), .Q(\mem[240][13] ) );
  DFQD1 \mem_reg[240][12]  ( .D(n825), .CP(clk), .Q(\mem[240][12] ) );
  DFQD1 \mem_reg[240][11]  ( .D(n824), .CP(clk), .Q(\mem[240][11] ) );
  DFQD1 \mem_reg[240][10]  ( .D(n823), .CP(clk), .Q(\mem[240][10] ) );
  DFQD1 \mem_reg[240][9]  ( .D(n822), .CP(clk), .Q(\mem[240][9] ) );
  DFQD1 \mem_reg[240][8]  ( .D(n821), .CP(clk), .Q(\mem[240][8] ) );
  DFQD1 \mem_reg[240][7]  ( .D(n820), .CP(clk), .Q(\mem[240][7] ) );
  DFQD1 \mem_reg[240][6]  ( .D(n819), .CP(clk), .Q(\mem[240][6] ) );
  DFQD1 \mem_reg[240][5]  ( .D(n818), .CP(clk), .Q(\mem[240][5] ) );
  DFQD1 \mem_reg[240][4]  ( .D(n817), .CP(clk), .Q(\mem[240][4] ) );
  DFQD1 \mem_reg[240][3]  ( .D(n816), .CP(clk), .Q(\mem[240][3] ) );
  DFQD1 \mem_reg[240][2]  ( .D(n815), .CP(clk), .Q(\mem[240][2] ) );
  DFQD1 \mem_reg[240][1]  ( .D(n814), .CP(clk), .Q(\mem[240][1] ) );
  DFQD1 \mem_reg[240][0]  ( .D(n813), .CP(clk), .Q(\mem[240][0] ) );
  DFQD1 \mem_reg[241][15]  ( .D(n812), .CP(clk), .Q(\mem[241][15] ) );
  DFQD1 \mem_reg[241][14]  ( .D(n811), .CP(clk), .Q(\mem[241][14] ) );
  DFQD1 \mem_reg[241][13]  ( .D(n810), .CP(clk), .Q(\mem[241][13] ) );
  DFQD1 \mem_reg[241][12]  ( .D(n809), .CP(clk), .Q(\mem[241][12] ) );
  DFQD1 \mem_reg[241][11]  ( .D(n808), .CP(clk), .Q(\mem[241][11] ) );
  DFQD1 \mem_reg[241][10]  ( .D(n807), .CP(clk), .Q(\mem[241][10] ) );
  DFQD1 \mem_reg[241][9]  ( .D(n806), .CP(clk), .Q(\mem[241][9] ) );
  DFQD1 \mem_reg[241][8]  ( .D(n805), .CP(clk), .Q(\mem[241][8] ) );
  DFQD1 \mem_reg[241][7]  ( .D(n804), .CP(clk), .Q(\mem[241][7] ) );
  DFQD1 \mem_reg[241][6]  ( .D(n803), .CP(clk), .Q(\mem[241][6] ) );
  DFQD1 \mem_reg[241][5]  ( .D(n802), .CP(clk), .Q(\mem[241][5] ) );
  DFQD1 \mem_reg[241][4]  ( .D(n801), .CP(clk), .Q(\mem[241][4] ) );
  DFQD1 \mem_reg[241][3]  ( .D(n800), .CP(clk), .Q(\mem[241][3] ) );
  DFQD1 \mem_reg[241][2]  ( .D(n799), .CP(clk), .Q(\mem[241][2] ) );
  DFQD1 \mem_reg[241][1]  ( .D(n798), .CP(clk), .Q(\mem[241][1] ) );
  DFQD1 \mem_reg[241][0]  ( .D(n797), .CP(clk), .Q(\mem[241][0] ) );
  DFQD1 \mem_reg[242][15]  ( .D(n796), .CP(clk), .Q(\mem[242][15] ) );
  DFQD1 \mem_reg[242][14]  ( .D(n795), .CP(clk), .Q(\mem[242][14] ) );
  DFQD1 \mem_reg[242][13]  ( .D(n794), .CP(clk), .Q(\mem[242][13] ) );
  DFQD1 \mem_reg[242][12]  ( .D(n793), .CP(clk), .Q(\mem[242][12] ) );
  DFQD1 \mem_reg[242][11]  ( .D(n792), .CP(clk), .Q(\mem[242][11] ) );
  DFQD1 \mem_reg[242][10]  ( .D(n791), .CP(clk), .Q(\mem[242][10] ) );
  DFQD1 \mem_reg[242][9]  ( .D(n790), .CP(clk), .Q(\mem[242][9] ) );
  DFQD1 \mem_reg[242][8]  ( .D(n789), .CP(clk), .Q(\mem[242][8] ) );
  DFQD1 \mem_reg[242][7]  ( .D(n788), .CP(clk), .Q(\mem[242][7] ) );
  DFQD1 \mem_reg[242][6]  ( .D(n787), .CP(clk), .Q(\mem[242][6] ) );
  DFQD1 \mem_reg[242][5]  ( .D(n786), .CP(clk), .Q(\mem[242][5] ) );
  DFQD1 \mem_reg[242][4]  ( .D(n785), .CP(clk), .Q(\mem[242][4] ) );
  DFQD1 \mem_reg[242][3]  ( .D(n784), .CP(clk), .Q(\mem[242][3] ) );
  DFQD1 \mem_reg[242][2]  ( .D(n783), .CP(clk), .Q(\mem[242][2] ) );
  DFQD1 \mem_reg[242][1]  ( .D(n782), .CP(clk), .Q(\mem[242][1] ) );
  DFQD1 \mem_reg[242][0]  ( .D(n781), .CP(clk), .Q(\mem[242][0] ) );
  DFQD1 \mem_reg[243][15]  ( .D(n780), .CP(clk), .Q(\mem[243][15] ) );
  DFQD1 \mem_reg[243][14]  ( .D(n779), .CP(clk), .Q(\mem[243][14] ) );
  DFQD1 \mem_reg[243][13]  ( .D(n778), .CP(clk), .Q(\mem[243][13] ) );
  DFQD1 \mem_reg[243][12]  ( .D(n777), .CP(clk), .Q(\mem[243][12] ) );
  DFQD1 \mem_reg[243][11]  ( .D(n776), .CP(clk), .Q(\mem[243][11] ) );
  DFQD1 \mem_reg[243][10]  ( .D(n775), .CP(clk), .Q(\mem[243][10] ) );
  DFQD1 \mem_reg[243][9]  ( .D(n774), .CP(clk), .Q(\mem[243][9] ) );
  DFQD1 \mem_reg[243][8]  ( .D(n773), .CP(clk), .Q(\mem[243][8] ) );
  DFQD1 \mem_reg[243][7]  ( .D(n772), .CP(clk), .Q(\mem[243][7] ) );
  DFQD1 \mem_reg[243][6]  ( .D(n771), .CP(clk), .Q(\mem[243][6] ) );
  DFQD1 \mem_reg[243][5]  ( .D(n770), .CP(clk), .Q(\mem[243][5] ) );
  DFQD1 \mem_reg[243][4]  ( .D(n769), .CP(clk), .Q(\mem[243][4] ) );
  DFQD1 \mem_reg[243][3]  ( .D(n768), .CP(clk), .Q(\mem[243][3] ) );
  DFQD1 \mem_reg[243][2]  ( .D(n767), .CP(clk), .Q(\mem[243][2] ) );
  DFQD1 \mem_reg[243][1]  ( .D(n766), .CP(clk), .Q(\mem[243][1] ) );
  DFQD1 \mem_reg[243][0]  ( .D(n765), .CP(clk), .Q(\mem[243][0] ) );
  DFQD1 \mem_reg[244][15]  ( .D(n764), .CP(clk), .Q(\mem[244][15] ) );
  DFQD1 \mem_reg[244][14]  ( .D(n763), .CP(clk), .Q(\mem[244][14] ) );
  DFQD1 \mem_reg[244][13]  ( .D(n762), .CP(clk), .Q(\mem[244][13] ) );
  DFQD1 \mem_reg[244][12]  ( .D(n761), .CP(clk), .Q(\mem[244][12] ) );
  DFQD1 \mem_reg[244][11]  ( .D(n760), .CP(clk), .Q(\mem[244][11] ) );
  DFQD1 \mem_reg[244][10]  ( .D(n759), .CP(clk), .Q(\mem[244][10] ) );
  DFQD1 \mem_reg[244][9]  ( .D(n758), .CP(clk), .Q(\mem[244][9] ) );
  DFQD1 \mem_reg[244][8]  ( .D(n757), .CP(clk), .Q(\mem[244][8] ) );
  DFQD1 \mem_reg[244][7]  ( .D(n756), .CP(clk), .Q(\mem[244][7] ) );
  DFQD1 \mem_reg[244][6]  ( .D(n755), .CP(clk), .Q(\mem[244][6] ) );
  DFQD1 \mem_reg[244][5]  ( .D(n754), .CP(clk), .Q(\mem[244][5] ) );
  DFQD1 \mem_reg[244][4]  ( .D(n753), .CP(clk), .Q(\mem[244][4] ) );
  DFQD1 \mem_reg[244][3]  ( .D(n752), .CP(clk), .Q(\mem[244][3] ) );
  DFQD1 \mem_reg[244][2]  ( .D(n751), .CP(clk), .Q(\mem[244][2] ) );
  DFQD1 \mem_reg[244][1]  ( .D(n750), .CP(clk), .Q(\mem[244][1] ) );
  DFQD1 \mem_reg[244][0]  ( .D(n749), .CP(clk), .Q(\mem[244][0] ) );
  DFQD1 \mem_reg[245][15]  ( .D(n748), .CP(clk), .Q(\mem[245][15] ) );
  DFQD1 \mem_reg[245][14]  ( .D(n747), .CP(clk), .Q(\mem[245][14] ) );
  DFQD1 \mem_reg[245][13]  ( .D(n746), .CP(clk), .Q(\mem[245][13] ) );
  DFQD1 \mem_reg[245][12]  ( .D(n745), .CP(clk), .Q(\mem[245][12] ) );
  DFQD1 \mem_reg[245][11]  ( .D(n744), .CP(clk), .Q(\mem[245][11] ) );
  DFQD1 \mem_reg[245][10]  ( .D(n743), .CP(clk), .Q(\mem[245][10] ) );
  DFQD1 \mem_reg[245][9]  ( .D(n742), .CP(clk), .Q(\mem[245][9] ) );
  DFQD1 \mem_reg[245][8]  ( .D(n741), .CP(clk), .Q(\mem[245][8] ) );
  DFQD1 \mem_reg[245][7]  ( .D(n740), .CP(clk), .Q(\mem[245][7] ) );
  DFQD1 \mem_reg[245][6]  ( .D(n739), .CP(clk), .Q(\mem[245][6] ) );
  DFQD1 \mem_reg[245][5]  ( .D(n738), .CP(clk), .Q(\mem[245][5] ) );
  DFQD1 \mem_reg[245][4]  ( .D(n737), .CP(clk), .Q(\mem[245][4] ) );
  DFQD1 \mem_reg[245][3]  ( .D(n736), .CP(clk), .Q(\mem[245][3] ) );
  DFQD1 \mem_reg[245][2]  ( .D(n735), .CP(clk), .Q(\mem[245][2] ) );
  DFQD1 \mem_reg[245][1]  ( .D(n734), .CP(clk), .Q(\mem[245][1] ) );
  DFQD1 \mem_reg[245][0]  ( .D(n733), .CP(clk), .Q(\mem[245][0] ) );
  DFQD1 \mem_reg[246][15]  ( .D(n732), .CP(clk), .Q(\mem[246][15] ) );
  DFQD1 \mem_reg[246][14]  ( .D(n731), .CP(clk), .Q(\mem[246][14] ) );
  DFQD1 \mem_reg[246][13]  ( .D(n730), .CP(clk), .Q(\mem[246][13] ) );
  DFQD1 \mem_reg[246][12]  ( .D(n729), .CP(clk), .Q(\mem[246][12] ) );
  DFQD1 \mem_reg[246][11]  ( .D(n728), .CP(clk), .Q(\mem[246][11] ) );
  DFQD1 \mem_reg[246][10]  ( .D(n727), .CP(clk), .Q(\mem[246][10] ) );
  DFQD1 \mem_reg[246][9]  ( .D(n726), .CP(clk), .Q(\mem[246][9] ) );
  DFQD1 \mem_reg[246][8]  ( .D(n725), .CP(clk), .Q(\mem[246][8] ) );
  DFQD1 \mem_reg[246][7]  ( .D(n724), .CP(clk), .Q(\mem[246][7] ) );
  DFQD1 \mem_reg[246][6]  ( .D(n723), .CP(clk), .Q(\mem[246][6] ) );
  DFQD1 \mem_reg[246][5]  ( .D(n722), .CP(clk), .Q(\mem[246][5] ) );
  DFQD1 \mem_reg[246][4]  ( .D(n721), .CP(clk), .Q(\mem[246][4] ) );
  DFQD1 \mem_reg[246][3]  ( .D(n720), .CP(clk), .Q(\mem[246][3] ) );
  DFQD1 \mem_reg[246][2]  ( .D(n719), .CP(clk), .Q(\mem[246][2] ) );
  DFQD1 \mem_reg[246][1]  ( .D(n718), .CP(clk), .Q(\mem[246][1] ) );
  DFQD1 \mem_reg[246][0]  ( .D(n717), .CP(clk), .Q(\mem[246][0] ) );
  DFQD1 \mem_reg[247][15]  ( .D(n716), .CP(clk), .Q(\mem[247][15] ) );
  DFQD1 \mem_reg[247][14]  ( .D(n715), .CP(clk), .Q(\mem[247][14] ) );
  DFQD1 \mem_reg[247][13]  ( .D(n714), .CP(clk), .Q(\mem[247][13] ) );
  DFQD1 \mem_reg[247][12]  ( .D(n713), .CP(clk), .Q(\mem[247][12] ) );
  DFQD1 \mem_reg[247][11]  ( .D(n712), .CP(clk), .Q(\mem[247][11] ) );
  DFQD1 \mem_reg[247][10]  ( .D(n711), .CP(clk), .Q(\mem[247][10] ) );
  DFQD1 \mem_reg[247][9]  ( .D(n710), .CP(clk), .Q(\mem[247][9] ) );
  DFQD1 \mem_reg[247][8]  ( .D(n709), .CP(clk), .Q(\mem[247][8] ) );
  DFQD1 \mem_reg[247][7]  ( .D(n708), .CP(clk), .Q(\mem[247][7] ) );
  DFQD1 \mem_reg[247][6]  ( .D(n707), .CP(clk), .Q(\mem[247][6] ) );
  DFQD1 \mem_reg[247][5]  ( .D(n706), .CP(clk), .Q(\mem[247][5] ) );
  DFQD1 \mem_reg[247][4]  ( .D(n705), .CP(clk), .Q(\mem[247][4] ) );
  DFQD1 \mem_reg[247][3]  ( .D(n704), .CP(clk), .Q(\mem[247][3] ) );
  DFQD1 \mem_reg[247][2]  ( .D(n703), .CP(clk), .Q(\mem[247][2] ) );
  DFQD1 \mem_reg[247][1]  ( .D(n702), .CP(clk), .Q(\mem[247][1] ) );
  DFQD1 \mem_reg[247][0]  ( .D(n701), .CP(clk), .Q(\mem[247][0] ) );
  DFQD1 \mem_reg[248][15]  ( .D(n700), .CP(clk), .Q(\mem[248][15] ) );
  DFQD1 \mem_reg[248][14]  ( .D(n699), .CP(clk), .Q(\mem[248][14] ) );
  DFQD1 \mem_reg[248][13]  ( .D(n698), .CP(clk), .Q(\mem[248][13] ) );
  DFQD1 \mem_reg[248][12]  ( .D(n697), .CP(clk), .Q(\mem[248][12] ) );
  DFQD1 \mem_reg[248][11]  ( .D(n696), .CP(clk), .Q(\mem[248][11] ) );
  DFQD1 \mem_reg[248][10]  ( .D(n695), .CP(clk), .Q(\mem[248][10] ) );
  DFQD1 \mem_reg[248][9]  ( .D(n694), .CP(clk), .Q(\mem[248][9] ) );
  DFQD1 \mem_reg[248][8]  ( .D(n693), .CP(clk), .Q(\mem[248][8] ) );
  DFQD1 \mem_reg[248][7]  ( .D(n692), .CP(clk), .Q(\mem[248][7] ) );
  DFQD1 \mem_reg[248][6]  ( .D(n691), .CP(clk), .Q(\mem[248][6] ) );
  DFQD1 \mem_reg[248][5]  ( .D(n690), .CP(clk), .Q(\mem[248][5] ) );
  DFQD1 \mem_reg[248][4]  ( .D(n689), .CP(clk), .Q(\mem[248][4] ) );
  DFQD1 \mem_reg[248][3]  ( .D(n688), .CP(clk), .Q(\mem[248][3] ) );
  DFQD1 \mem_reg[248][2]  ( .D(n687), .CP(clk), .Q(\mem[248][2] ) );
  DFQD1 \mem_reg[248][1]  ( .D(n686), .CP(clk), .Q(\mem[248][1] ) );
  DFQD1 \mem_reg[248][0]  ( .D(n685), .CP(clk), .Q(\mem[248][0] ) );
  DFQD1 \mem_reg[249][15]  ( .D(n684), .CP(clk), .Q(\mem[249][15] ) );
  DFQD1 \mem_reg[249][14]  ( .D(n683), .CP(clk), .Q(\mem[249][14] ) );
  DFQD1 \mem_reg[249][13]  ( .D(n682), .CP(clk), .Q(\mem[249][13] ) );
  DFQD1 \mem_reg[249][12]  ( .D(n681), .CP(clk), .Q(\mem[249][12] ) );
  DFQD1 \mem_reg[249][11]  ( .D(n680), .CP(clk), .Q(\mem[249][11] ) );
  DFQD1 \mem_reg[249][10]  ( .D(n679), .CP(clk), .Q(\mem[249][10] ) );
  DFQD1 \mem_reg[249][9]  ( .D(n678), .CP(clk), .Q(\mem[249][9] ) );
  DFQD1 \mem_reg[249][8]  ( .D(n677), .CP(clk), .Q(\mem[249][8] ) );
  DFQD1 \mem_reg[249][7]  ( .D(n676), .CP(clk), .Q(\mem[249][7] ) );
  DFQD1 \mem_reg[249][6]  ( .D(n675), .CP(clk), .Q(\mem[249][6] ) );
  DFQD1 \mem_reg[249][5]  ( .D(n674), .CP(clk), .Q(\mem[249][5] ) );
  DFQD1 \mem_reg[249][4]  ( .D(n673), .CP(clk), .Q(\mem[249][4] ) );
  DFQD1 \mem_reg[249][3]  ( .D(n672), .CP(clk), .Q(\mem[249][3] ) );
  DFQD1 \mem_reg[249][2]  ( .D(n671), .CP(clk), .Q(\mem[249][2] ) );
  DFQD1 \mem_reg[249][1]  ( .D(n670), .CP(clk), .Q(\mem[249][1] ) );
  DFQD1 \mem_reg[249][0]  ( .D(n669), .CP(clk), .Q(\mem[249][0] ) );
  DFQD1 \mem_reg[250][15]  ( .D(n668), .CP(clk), .Q(\mem[250][15] ) );
  DFQD1 \mem_reg[250][14]  ( .D(n667), .CP(clk), .Q(\mem[250][14] ) );
  DFQD1 \mem_reg[250][13]  ( .D(n666), .CP(clk), .Q(\mem[250][13] ) );
  DFQD1 \mem_reg[250][12]  ( .D(n665), .CP(clk), .Q(\mem[250][12] ) );
  DFQD1 \mem_reg[250][11]  ( .D(n664), .CP(clk), .Q(\mem[250][11] ) );
  DFQD1 \mem_reg[250][10]  ( .D(n663), .CP(clk), .Q(\mem[250][10] ) );
  DFQD1 \mem_reg[250][9]  ( .D(n662), .CP(clk), .Q(\mem[250][9] ) );
  DFQD1 \mem_reg[250][8]  ( .D(n661), .CP(clk), .Q(\mem[250][8] ) );
  DFQD1 \mem_reg[250][7]  ( .D(n660), .CP(clk), .Q(\mem[250][7] ) );
  DFQD1 \mem_reg[250][6]  ( .D(n659), .CP(clk), .Q(\mem[250][6] ) );
  DFQD1 \mem_reg[250][5]  ( .D(n658), .CP(clk), .Q(\mem[250][5] ) );
  DFQD1 \mem_reg[250][4]  ( .D(n657), .CP(clk), .Q(\mem[250][4] ) );
  DFQD1 \mem_reg[250][3]  ( .D(n656), .CP(clk), .Q(\mem[250][3] ) );
  DFQD1 \mem_reg[250][2]  ( .D(n655), .CP(clk), .Q(\mem[250][2] ) );
  DFQD1 \mem_reg[250][1]  ( .D(n654), .CP(clk), .Q(\mem[250][1] ) );
  DFQD1 \mem_reg[250][0]  ( .D(n653), .CP(clk), .Q(\mem[250][0] ) );
  DFQD1 \mem_reg[251][15]  ( .D(n652), .CP(clk), .Q(\mem[251][15] ) );
  DFQD1 \mem_reg[251][14]  ( .D(n651), .CP(clk), .Q(\mem[251][14] ) );
  DFQD1 \mem_reg[251][13]  ( .D(n650), .CP(clk), .Q(\mem[251][13] ) );
  DFQD1 \mem_reg[251][12]  ( .D(n649), .CP(clk), .Q(\mem[251][12] ) );
  DFQD1 \mem_reg[251][11]  ( .D(n648), .CP(clk), .Q(\mem[251][11] ) );
  DFQD1 \mem_reg[251][10]  ( .D(n647), .CP(clk), .Q(\mem[251][10] ) );
  DFQD1 \mem_reg[251][9]  ( .D(n646), .CP(clk), .Q(\mem[251][9] ) );
  DFQD1 \mem_reg[251][8]  ( .D(n645), .CP(clk), .Q(\mem[251][8] ) );
  DFQD1 \mem_reg[251][7]  ( .D(n644), .CP(clk), .Q(\mem[251][7] ) );
  DFQD1 \mem_reg[251][6]  ( .D(n643), .CP(clk), .Q(\mem[251][6] ) );
  DFQD1 \mem_reg[251][5]  ( .D(n642), .CP(clk), .Q(\mem[251][5] ) );
  DFQD1 \mem_reg[251][4]  ( .D(n641), .CP(clk), .Q(\mem[251][4] ) );
  DFQD1 \mem_reg[251][3]  ( .D(n640), .CP(clk), .Q(\mem[251][3] ) );
  DFQD1 \mem_reg[251][2]  ( .D(n639), .CP(clk), .Q(\mem[251][2] ) );
  DFQD1 \mem_reg[251][1]  ( .D(n638), .CP(clk), .Q(\mem[251][1] ) );
  DFQD1 \mem_reg[251][0]  ( .D(n637), .CP(clk), .Q(\mem[251][0] ) );
  DFQD1 \mem_reg[252][15]  ( .D(n636), .CP(clk), .Q(\mem[252][15] ) );
  DFQD1 \mem_reg[252][14]  ( .D(n635), .CP(clk), .Q(\mem[252][14] ) );
  DFQD1 \mem_reg[252][13]  ( .D(n634), .CP(clk), .Q(\mem[252][13] ) );
  DFQD1 \mem_reg[252][12]  ( .D(n633), .CP(clk), .Q(\mem[252][12] ) );
  DFQD1 \mem_reg[252][11]  ( .D(n632), .CP(clk), .Q(\mem[252][11] ) );
  DFQD1 \mem_reg[252][10]  ( .D(n631), .CP(clk), .Q(\mem[252][10] ) );
  DFQD1 \mem_reg[252][9]  ( .D(n630), .CP(clk), .Q(\mem[252][9] ) );
  DFQD1 \mem_reg[252][8]  ( .D(n629), .CP(clk), .Q(\mem[252][8] ) );
  DFQD1 \mem_reg[252][7]  ( .D(n628), .CP(clk), .Q(\mem[252][7] ) );
  DFQD1 \mem_reg[252][6]  ( .D(n627), .CP(clk), .Q(\mem[252][6] ) );
  DFQD1 \mem_reg[252][5]  ( .D(n626), .CP(clk), .Q(\mem[252][5] ) );
  DFQD1 \mem_reg[252][4]  ( .D(n625), .CP(clk), .Q(\mem[252][4] ) );
  DFQD1 \mem_reg[252][3]  ( .D(n624), .CP(clk), .Q(\mem[252][3] ) );
  DFQD1 \mem_reg[252][2]  ( .D(n623), .CP(clk), .Q(\mem[252][2] ) );
  DFQD1 \mem_reg[252][1]  ( .D(n622), .CP(clk), .Q(\mem[252][1] ) );
  DFQD1 \mem_reg[252][0]  ( .D(n621), .CP(clk), .Q(\mem[252][0] ) );
  DFQD1 \mem_reg[253][15]  ( .D(n620), .CP(clk), .Q(\mem[253][15] ) );
  DFQD1 \mem_reg[253][14]  ( .D(n619), .CP(clk), .Q(\mem[253][14] ) );
  DFQD1 \mem_reg[253][13]  ( .D(n618), .CP(clk), .Q(\mem[253][13] ) );
  DFQD1 \mem_reg[253][12]  ( .D(n617), .CP(clk), .Q(\mem[253][12] ) );
  DFQD1 \mem_reg[253][11]  ( .D(n616), .CP(clk), .Q(\mem[253][11] ) );
  DFQD1 \mem_reg[253][10]  ( .D(n615), .CP(clk), .Q(\mem[253][10] ) );
  DFQD1 \mem_reg[253][9]  ( .D(n614), .CP(clk), .Q(\mem[253][9] ) );
  DFQD1 \mem_reg[253][8]  ( .D(n613), .CP(clk), .Q(\mem[253][8] ) );
  DFQD1 \mem_reg[253][7]  ( .D(n612), .CP(clk), .Q(\mem[253][7] ) );
  DFQD1 \mem_reg[253][6]  ( .D(n611), .CP(clk), .Q(\mem[253][6] ) );
  DFQD1 \mem_reg[253][5]  ( .D(n610), .CP(clk), .Q(\mem[253][5] ) );
  DFQD1 \mem_reg[253][4]  ( .D(n609), .CP(clk), .Q(\mem[253][4] ) );
  DFQD1 \mem_reg[253][3]  ( .D(n608), .CP(clk), .Q(\mem[253][3] ) );
  DFQD1 \mem_reg[253][2]  ( .D(n607), .CP(clk), .Q(\mem[253][2] ) );
  DFQD1 \mem_reg[253][1]  ( .D(n606), .CP(clk), .Q(\mem[253][1] ) );
  DFQD1 \mem_reg[253][0]  ( .D(n605), .CP(clk), .Q(\mem[253][0] ) );
  DFQD1 \mem_reg[254][15]  ( .D(n604), .CP(clk), .Q(\mem[254][15] ) );
  DFQD1 \mem_reg[254][14]  ( .D(n603), .CP(clk), .Q(\mem[254][14] ) );
  DFQD1 \mem_reg[254][13]  ( .D(n602), .CP(clk), .Q(\mem[254][13] ) );
  DFQD1 \mem_reg[254][12]  ( .D(n601), .CP(clk), .Q(\mem[254][12] ) );
  DFQD1 \mem_reg[254][11]  ( .D(n600), .CP(clk), .Q(\mem[254][11] ) );
  DFQD1 \mem_reg[254][10]  ( .D(n599), .CP(clk), .Q(\mem[254][10] ) );
  DFQD1 \mem_reg[254][9]  ( .D(n598), .CP(clk), .Q(\mem[254][9] ) );
  DFQD1 \mem_reg[254][8]  ( .D(n597), .CP(clk), .Q(\mem[254][8] ) );
  DFQD1 \mem_reg[254][7]  ( .D(n596), .CP(clk), .Q(\mem[254][7] ) );
  DFQD1 \mem_reg[254][6]  ( .D(n595), .CP(clk), .Q(\mem[254][6] ) );
  DFQD1 \mem_reg[254][5]  ( .D(n594), .CP(clk), .Q(\mem[254][5] ) );
  DFQD1 \mem_reg[254][4]  ( .D(n593), .CP(clk), .Q(\mem[254][4] ) );
  DFQD1 \mem_reg[254][3]  ( .D(n592), .CP(clk), .Q(\mem[254][3] ) );
  DFQD1 \mem_reg[254][2]  ( .D(n591), .CP(clk), .Q(\mem[254][2] ) );
  DFQD1 \mem_reg[254][1]  ( .D(n590), .CP(clk), .Q(\mem[254][1] ) );
  DFQD1 \mem_reg[254][0]  ( .D(n589), .CP(clk), .Q(\mem[254][0] ) );
  DFQD1 \mem_reg[255][15]  ( .D(n588), .CP(clk), .Q(\mem[255][15] ) );
  DFQD1 \mem_reg[255][14]  ( .D(n587), .CP(clk), .Q(\mem[255][14] ) );
  DFQD1 \mem_reg[255][13]  ( .D(n586), .CP(clk), .Q(\mem[255][13] ) );
  DFQD1 \mem_reg[255][12]  ( .D(n585), .CP(clk), .Q(\mem[255][12] ) );
  DFQD1 \mem_reg[255][11]  ( .D(n584), .CP(clk), .Q(\mem[255][11] ) );
  DFQD1 \mem_reg[255][10]  ( .D(n583), .CP(clk), .Q(\mem[255][10] ) );
  DFQD1 \mem_reg[255][9]  ( .D(n582), .CP(clk), .Q(\mem[255][9] ) );
  DFQD1 \mem_reg[255][8]  ( .D(n581), .CP(clk), .Q(\mem[255][8] ) );
  DFQD1 \mem_reg[255][7]  ( .D(n580), .CP(clk), .Q(\mem[255][7] ) );
  DFQD1 \mem_reg[255][6]  ( .D(n579), .CP(clk), .Q(\mem[255][6] ) );
  DFQD1 \mem_reg[255][5]  ( .D(n578), .CP(clk), .Q(\mem[255][5] ) );
  DFQD1 \mem_reg[255][4]  ( .D(n577), .CP(clk), .Q(\mem[255][4] ) );
  DFQD1 \mem_reg[255][3]  ( .D(n576), .CP(clk), .Q(\mem[255][3] ) );
  DFQD1 \mem_reg[255][2]  ( .D(n575), .CP(clk), .Q(\mem[255][2] ) );
  DFQD1 \mem_reg[255][1]  ( .D(n574), .CP(clk), .Q(\mem[255][1] ) );
  DFQD1 \mem_reg[255][0]  ( .D(n573), .CP(clk), .Q(\mem[255][0] ) );
  NR2D0 U2 ( .A1(n71), .A2(n53), .ZN(n5966) );
  AOI22D0 U3 ( .A1(n6759), .A2(\mem[206][12] ), .B1(n6809), .B2(\mem[201][12] ), .ZN(n5116) );
  AOI22D0 U4 ( .A1(n6953), .A2(\mem[239][12] ), .B1(n6988), .B2(\mem[255][12] ), .ZN(n5095) );
  AOI22D0 U5 ( .A1(n6179), .A2(\mem[111][12] ), .B1(n6760), .B2(\mem[109][12] ), .ZN(n5072) );
  AOI22D0 U6 ( .A1(n6830), .A2(\mem[71][12] ), .B1(n6891), .B2(\mem[90][12] ), 
        .ZN(n5059) );
  AOI22D0 U7 ( .A1(n6881), .A2(\mem[144][12] ), .B1(n6923), .B2(\mem[162][12] ), .ZN(n5036) );
  AOI22D0 U8 ( .A1(n6913), .A2(\mem[155][12] ), .B1(n6993), .B2(\mem[181][12] ), .ZN(n5015) );
  AOI22D0 U9 ( .A1(n6892), .A2(\mem[44][15] ), .B1(n6923), .B2(\mem[34][15] ), 
        .ZN(n4764) );
  AOI22D0 U10 ( .A1(n6981), .A2(\mem[60][15] ), .B1(n6905), .B2(\mem[59][15] ), 
        .ZN(n4743) );
  AOI22D0 U11 ( .A1(n6994), .A2(\mem[254][15] ), .B1(n6871), .B2(
        \mem[249][15] ), .ZN(n4720) );
  AOI22D0 U12 ( .A1(n6991), .A2(\mem[212][15] ), .B1(n6906), .B2(
        \mem[204][15] ), .ZN(n4707) );
  AOI22D0 U13 ( .A1(n6747), .A2(\mem[84][15] ), .B1(n6728), .B2(\mem[116][15] ), .ZN(n4684) );
  AOI22D0 U14 ( .A1(n6530), .A2(\mem[123][15] ), .B1(n6874), .B2(
        \mem[106][15] ), .ZN(n567) );
  AOI22D0 U15 ( .A1(n6859), .A2(\mem[52][14] ), .B1(n6965), .B2(\mem[13][14] ), 
        .ZN(n4938) );
  AOI22D0 U16 ( .A1(n6966), .A2(\mem[50][14] ), .B1(n6748), .B2(\mem[41][14] ), 
        .ZN(n4925) );
  AOI22D0 U17 ( .A1(n6165), .A2(\mem[238][14] ), .B1(n6966), .B2(
        \mem[242][14] ), .ZN(n4902) );
  AOI22D0 U18 ( .A1(n6969), .A2(\mem[210][14] ), .B1(n6888), .B2(
        \mem[192][14] ), .ZN(n4881) );
  AOI22D0 U19 ( .A1(n6905), .A2(\mem[187][14] ), .B1(n6957), .B2(
        \mem[185][14] ), .ZN(n4858) );
  AOI22D0 U20 ( .A1(n6747), .A2(\mem[148][14] ), .B1(n6748), .B2(
        \mem[169][14] ), .ZN(n4845) );
  AOI22D0 U21 ( .A1(n6979), .A2(\mem[78][11] ), .B1(n6707), .B2(\mem[87][11] ), 
        .ZN(n5290) );
  AOI22D0 U22 ( .A1(n6525), .A2(\mem[99][11] ), .B1(n6883), .B2(\mem[112][11] ), .ZN(n5281) );
  AOI22D0 U23 ( .A1(n6872), .A2(\mem[70][11] ), .B1(n6926), .B2(\mem[65][11] ), 
        .ZN(n5260) );
  AOI22D0 U24 ( .A1(n6914), .A2(\mem[197][11] ), .B1(n6563), .B2(
        \mem[200][11] ), .ZN(n5237) );
  AOI22D0 U25 ( .A1(n6847), .A2(\mem[217][11] ), .B1(n6728), .B2(
        \mem[244][11] ), .ZN(n5216) );
  AOI22D0 U26 ( .A1(n6165), .A2(\mem[174][11] ), .B1(n6904), .B2(
        \mem[147][11] ), .ZN(n5201) );
  AOI22D0 U27 ( .A1(n6883), .A2(\mem[176][11] ), .B1(n6748), .B2(
        \mem[169][11] ), .ZN(n5180) );
  AOI22D0 U28 ( .A1(n6874), .A2(\mem[234][6] ), .B1(n6915), .B2(\mem[205][6] ), 
        .ZN(n6144) );
  AOI22D0 U29 ( .A1(n6863), .A2(\mem[247][6] ), .B1(n6988), .B2(\mem[255][6] ), 
        .ZN(n6123) );
  AOI22D0 U30 ( .A1(n6922), .A2(\mem[29][6] ), .B1(n6862), .B2(\mem[40][6] ), 
        .ZN(n6108) );
  AOI22D0 U31 ( .A1(n6959), .A2(\mem[3][6] ), .B1(n6968), .B2(\mem[41][6] ), 
        .ZN(n6087) );
  AOI22D0 U32 ( .A1(n6890), .A2(\mem[100][6] ), .B1(n6959), .B2(\mem[67][6] ), 
        .ZN(n6064) );
  AOI22D0 U33 ( .A1(n6754), .A2(\mem[69][6] ), .B1(n6563), .B2(\mem[72][6] ), 
        .ZN(n6043) );
  AOI22D0 U34 ( .A1(n6979), .A2(\mem[206][10] ), .B1(n6958), .B2(
        \mem[209][10] ), .ZN(n5809) );
  AOI22D0 U35 ( .A1(n6934), .A2(\mem[216][10] ), .B1(n6966), .B2(
        \mem[242][10] ), .ZN(n5788) );
  AOI22D0 U36 ( .A1(n6775), .A2(\mem[44][10] ), .B1(n6860), .B2(\mem[35][10] ), 
        .ZN(n5765) );
  AOI22D0 U37 ( .A1(n6991), .A2(\mem[20][10] ), .B1(n6916), .B2(\mem[21][10] ), 
        .ZN(n5744) );
  AOI22D0 U38 ( .A1(n6923), .A2(\mem[34][10] ), .B1(n6789), .B2(\mem[62][10] ), 
        .ZN(n5735) );
  AOI22D0 U39 ( .A1(n6924), .A2(\mem[160][10] ), .B1(n6837), .B2(
        \mem[143][10] ), .ZN(n5712) );
  AOI22D0 U40 ( .A1(n6971), .A2(\mem[166][10] ), .B1(n6904), .B2(
        \mem[147][10] ), .ZN(n5691) );
  AOI22D0 U41 ( .A1(n6773), .A2(\mem[228][9] ), .B1(n6928), .B2(\mem[199][9] ), 
        .ZN(n5967) );
  AOI22D0 U42 ( .A1(n6883), .A2(\mem[240][9] ), .B1(n6791), .B2(\mem[224][9] ), 
        .ZN(n5953) );
  AOI22D0 U43 ( .A1(n6923), .A2(\mem[34][9] ), .B1(n6847), .B2(\mem[25][9] ), 
        .ZN(n5930) );
  AOI22D0 U44 ( .A1(n6784), .A2(\mem[28][9] ), .B1(n6639), .B2(\mem[39][9] ), 
        .ZN(n5909) );
  AOI22D0 U45 ( .A1(n6803), .A2(\mem[119][9] ), .B1(n6174), .B2(\mem[118][9] ), 
        .ZN(n5886) );
  AOI22D0 U46 ( .A1(n6728), .A2(\mem[116][9] ), .B1(n6748), .B2(\mem[105][9] ), 
        .ZN(n5873) );
  AOI22D0 U47 ( .A1(n6980), .A2(\mem[125][8] ), .B1(n6903), .B2(\mem[115][8] ), 
        .ZN(n5632) );
  AOI22D0 U48 ( .A1(n6784), .A2(\mem[92][8] ), .B1(n6902), .B2(\mem[101][8] ), 
        .ZN(n5611) );
  AOI22D0 U49 ( .A1(n6790), .A2(\mem[219][8] ), .B1(n6174), .B2(\mem[246][8] ), 
        .ZN(n5588) );
  AOI22D0 U50 ( .A1(n6915), .A2(\mem[205][8] ), .B1(n6902), .B2(\mem[229][8] ), 
        .ZN(n5575) );
  AOI22D0 U51 ( .A1(n6957), .A2(\mem[185][8] ), .B1(n6978), .B2(\mem[136][8] ), 
        .ZN(n5552) );
  AOI22D0 U52 ( .A1(n6889), .A2(\mem[156][8] ), .B1(n6995), .B2(\mem[151][8] ), 
        .ZN(n5531) );
  AOI22D0 U53 ( .A1(n6904), .A2(\mem[211][7] ), .B1(n6915), .B2(\mem[205][7] ), 
        .ZN(n6330) );
  AOI22D0 U54 ( .A1(n6979), .A2(\mem[206][7] ), .B1(n6707), .B2(\mem[215][7] ), 
        .ZN(n6320) );
  AOI22D0 U55 ( .A1(n6890), .A2(\mem[228][7] ), .B1(n6889), .B2(\mem[220][7] ), 
        .ZN(n6299) );
  AOI22D0 U56 ( .A1(n6879), .A2(\mem[58][7] ), .B1(n6916), .B2(\mem[21][7] ), 
        .ZN(n6275) );
  AOI22D0 U57 ( .A1(n6639), .A2(\mem[39][7] ), .B1(n6698), .B2(\mem[2][7] ), 
        .ZN(n6254) );
  AOI22D0 U58 ( .A1(n6928), .A2(\mem[135][7] ), .B1(n6869), .B2(\mem[177][7] ), 
        .ZN(n6239) );
  AOI22D0 U59 ( .A1(n6863), .A2(\mem[183][7] ), .B1(n6748), .B2(\mem[169][7] ), 
        .ZN(n6218) );
  ND4D0 U60 ( .A1(n5075), .A2(n5074), .A3(n5073), .A4(n5072), .ZN(n5081) );
  AOI22D0 U61 ( .A1(n6448), .A2(\mem[192][13] ), .B1(n6906), .B2(
        \mem[204][13] ), .ZN(n504) );
  AOI22D0 U62 ( .A1(n6842), .A2(\mem[218][13] ), .B1(n6748), .B2(
        \mem[233][13] ), .ZN(n483) );
  AOI22D0 U63 ( .A1(n6914), .A2(\mem[5][13] ), .B1(n6774), .B2(\mem[49][13] ), 
        .ZN(n460) );
  AOI22D0 U64 ( .A1(n6847), .A2(\mem[25][13] ), .B1(n6936), .B2(\mem[17][13] ), 
        .ZN(n447) );
  AOI22D0 U65 ( .A1(n6953), .A2(\mem[175][13] ), .B1(n6890), .B2(
        \mem[164][13] ), .ZN(n424) );
  AOI22D0 U66 ( .A1(n6995), .A2(\mem[151][13] ), .B1(n6956), .B2(
        \mem[168][13] ), .ZN(n403) );
  ND4D0 U67 ( .A1(n4777), .A2(n4776), .A3(n4775), .A4(n4774), .ZN(n4778) );
  ND4D0 U68 ( .A1(n4703), .A2(n4702), .A3(n4701), .A4(n4700), .ZN(n4719) );
  ND4D0 U69 ( .A1(n4921), .A2(n4920), .A3(n4919), .A4(n4918), .ZN(n4932) );
  ND4D0 U70 ( .A1(n4841), .A2(n4840), .A3(n4839), .A4(n4838), .ZN(n4847) );
  ND4D0 U71 ( .A1(n5247), .A2(n5246), .A3(n5245), .A4(n5244), .ZN(n5253) );
  ND4D0 U72 ( .A1(n6154), .A2(n6153), .A3(n6152), .A4(n6151), .ZN(n6155) );
  ND4D0 U73 ( .A1(n6080), .A2(n6079), .A3(n6078), .A4(n6077), .ZN(n6096) );
  ND4D0 U74 ( .A1(n5781), .A2(n5780), .A3(n5779), .A4(n5778), .ZN(n5792) );
  ND4D0 U75 ( .A1(n5701), .A2(n5700), .A3(n5699), .A4(n5698), .ZN(n5707) );
  ND4D0 U76 ( .A1(n5919), .A2(n5918), .A3(n5917), .A4(n5916), .ZN(n5920) );
  ND4D0 U77 ( .A1(n5625), .A2(n5624), .A3(n5623), .A4(n5622), .ZN(n5641) );
  ND4D0 U78 ( .A1(n5545), .A2(n5544), .A3(n5543), .A4(n5542), .ZN(n5556) );
  ND4D0 U79 ( .A1(n6285), .A2(n6284), .A3(n6283), .A4(n6282), .ZN(n6291) );
  AOI22D0 U80 ( .A1(n6658), .A2(\mem[50][12] ), .B1(n6882), .B2(\mem[15][12] ), 
        .ZN(n5143) );
  AOI22D0 U81 ( .A1(n6530), .A2(\mem[59][12] ), .B1(n6728), .B2(\mem[52][12] ), 
        .ZN(n5134) );
  AOI22D0 U82 ( .A1(n6917), .A2(\mem[46][12] ), .B1(n6789), .B2(\mem[62][12] ), 
        .ZN(n4986) );
  AOI22D0 U83 ( .A1(n6748), .A2(\mem[233][4] ), .B1(n6915), .B2(\mem[205][4] ), 
        .ZN(n161) );
  AOI22D0 U84 ( .A1(n6728), .A2(\mem[244][4] ), .B1(n6760), .B2(\mem[237][4] ), 
        .ZN(n140) );
  AOI22D0 U85 ( .A1(n6959), .A2(\mem[67][4] ), .B1(n6837), .B2(\mem[79][4] ), 
        .ZN(n116) );
  AOI22D0 U86 ( .A1(n6995), .A2(\mem[87][4] ), .B1(n6738), .B2(\mem[101][4] ), 
        .ZN(n95) );
  AOI22D0 U87 ( .A1(n6970), .A2(\mem[144][4] ), .B1(n6879), .B2(\mem[186][4] ), 
        .ZN(n80) );
  AOI22D0 U88 ( .A1(n6888), .A2(\mem[128][4] ), .B1(n6774), .B2(\mem[177][4] ), 
        .ZN(n43) );
  ND4D0 U89 ( .A1(n505), .A2(n504), .A3(n503), .A4(n502), .ZN(n511) );
  ND4D0 U90 ( .A1(n425), .A2(n424), .A3(n423), .A4(n422), .ZN(n426) );
  AOI22D0 U91 ( .A1(n6969), .A2(\mem[146][15] ), .B1(n6881), .B2(
        \mem[144][15] ), .ZN(n4797) );
  AOI22D0 U92 ( .A1(n6871), .A2(\mem[185][15] ), .B1(n6862), .B2(
        \mem[168][15] ), .ZN(n554) );
  AOI22D0 U93 ( .A1(n6924), .A2(\mem[160][15] ), .B1(n6955), .B2(
        \mem[149][15] ), .ZN(n544) );
  AOI22D0 U94 ( .A1(n6892), .A2(\mem[108][14] ), .B1(n6993), .B2(
        \mem[117][14] ), .ZN(n4960) );
  AOI22D0 U95 ( .A1(n6890), .A2(\mem[100][14] ), .B1(n6905), .B2(
        \mem[123][14] ), .ZN(n4820) );
  AOI22D0 U96 ( .A1(n6967), .A2(\mem[231][2] ), .B1(n6988), .B2(\mem[255][2] ), 
        .ZN(n6492) );
  AOI22D0 U97 ( .A1(n6747), .A2(\mem[212][2] ), .B1(n6922), .B2(\mem[221][2] ), 
        .ZN(n6478) );
  AOI22D0 U98 ( .A1(n6989), .A2(\mem[70][2] ), .B1(n6933), .B2(\mem[97][2] ), 
        .ZN(n6455) );
  AOI22D0 U99 ( .A1(n6890), .A2(\mem[100][2] ), .B1(n6828), .B2(\mem[120][2] ), 
        .ZN(n6433) );
  AOI22D0 U100 ( .A1(n6891), .A2(\mem[154][2] ), .B1(n6936), .B2(\mem[145][2] ), .ZN(n6410) );
  AOI22D0 U101 ( .A1(n6971), .A2(\mem[166][2] ), .B1(n6966), .B2(\mem[178][2] ), .ZN(n6397) );
  AOI22D0 U102 ( .A1(n6773), .A2(\mem[228][3] ), .B1(n6925), .B2(\mem[237][3] ), .ZN(n6683) );
  AOI22D0 U103 ( .A1(n6860), .A2(\mem[227][3] ), .B1(n6789), .B2(\mem[254][3] ), .ZN(n6661) );
  AOI22D0 U104 ( .A1(n6927), .A2(\mem[25][3] ), .B1(n6774), .B2(\mem[49][3] ), 
        .ZN(n6635) );
  AOI22D0 U105 ( .A1(n6889), .A2(\mem[28][3] ), .B1(n6982), .B2(\mem[2][3] ), 
        .ZN(n6622) );
  AOI22D0 U106 ( .A1(n6917), .A2(\mem[174][3] ), .B1(n6880), .B2(\mem[139][3] ), .ZN(n6598) );
  AOI22D0 U107 ( .A1(n6913), .A2(\mem[155][3] ), .B1(n6906), .B2(\mem[140][3] ), .ZN(n6577) );
  AOI22D0 U108 ( .A1(n6983), .A2(\mem[48][11] ), .B1(n6837), .B2(\mem[15][11] ), .ZN(n5308) );
  AOI22D0 U109 ( .A1(n6923), .A2(\mem[34][11] ), .B1(n6774), .B2(\mem[49][11] ), .ZN(n5168) );
  AOI22D0 U110 ( .A1(n6862), .A2(\mem[168][6] ), .B1(n6978), .B2(\mem[136][6] ), .ZN(n6181) );
  AOI22D0 U111 ( .A1(n6861), .A2(\mem[132][6] ), .B1(n6936), .B2(\mem[145][6] ), .ZN(n6027) );
  AOI22D0 U112 ( .A1(n6892), .A2(\mem[172][6] ), .B1(n6955), .B2(\mem[149][6] ), .ZN(n6020) );
  AOI22D0 U113 ( .A1(n6809), .A2(\mem[73][10] ), .B1(n6922), .B2(\mem[93][10] ), .ZN(n5823) );
  AOI22D0 U114 ( .A1(n6525), .A2(\mem[99][10] ), .B1(n6971), .B2(
        \mem[102][10] ), .ZN(n5683) );
  AOI22D0 U115 ( .A1(n6883), .A2(\mem[176][9] ), .B1(n6923), .B2(\mem[162][9] ), .ZN(n6004) );
  AOI22D0 U116 ( .A1(n6914), .A2(\mem[133][9] ), .B1(n6658), .B2(\mem[178][9] ), .ZN(n5995) );
  AOI22D0 U117 ( .A1(n6913), .A2(\mem[155][9] ), .B1(n6924), .B2(\mem[160][9] ), .ZN(n5846) );
  AOI22D0 U118 ( .A1(n6829), .A2(\mem[38][8] ), .B1(n6680), .B2(\mem[31][8] ), 
        .ZN(n5658) );
  AOI22D0 U119 ( .A1(n6934), .A2(\mem[24][8] ), .B1(n6728), .B2(\mem[52][8] ), 
        .ZN(n5510) );
  AOI22D0 U120 ( .A1(n6970), .A2(\mem[16][8] ), .B1(n6804), .B2(\mem[19][8] ), 
        .ZN(n5501) );
  AOI22D0 U121 ( .A1(n6914), .A2(\mem[69][7] ), .B1(n6748), .B2(\mem[105][7] ), 
        .ZN(n6345) );
  AOI22D0 U122 ( .A1(n6749), .A2(\mem[107][7] ), .B1(n6925), .B2(\mem[109][7] ), .ZN(n6203) );
  CKND2D0 U123 ( .A1(n5043), .A2(n5042), .ZN(n5130) );
  ND4D0 U124 ( .A1(n118), .A2(n117), .A3(n116), .A4(n115), .ZN(n124) );
  AOI22D0 U125 ( .A1(n6934), .A2(\mem[216][5] ), .B1(n6928), .B2(\mem[199][5] ), .ZN(n5462) );
  AOI22D0 U126 ( .A1(n6179), .A2(\mem[239][5] ), .B1(n6869), .B2(\mem[241][5] ), .ZN(n5453) );
  AOI22D0 U127 ( .A1(n6325), .A2(\mem[203][5] ), .B1(n6847), .B2(\mem[217][5] ), .ZN(n5432) );
  AOI22D0 U128 ( .A1(n6971), .A2(\mem[102][5] ), .B1(n6873), .B2(\mem[94][5] ), 
        .ZN(n5409) );
  AOI22D0 U129 ( .A1(n6165), .A2(\mem[110][5] ), .B1(n6791), .B2(\mem[96][5] ), 
        .ZN(n5388) );
  AOI22D0 U130 ( .A1(n6754), .A2(\mem[133][5] ), .B1(n6563), .B2(\mem[136][5] ), .ZN(n5373) );
  AOI22D0 U131 ( .A1(n6804), .A2(\mem[147][5] ), .B1(n6965), .B2(\mem[141][5] ), .ZN(n5352) );
  AOI22D0 U132 ( .A1(n6803), .A2(\mem[119][13] ), .B1(n6658), .B2(
        \mem[114][13] ), .ZN(n523) );
  AOI22D0 U133 ( .A1(n6889), .A2(\mem[92][13] ), .B1(n6922), .B2(\mem[93][13] ), .ZN(n383) );
  ND4D0 U134 ( .A1(n4802), .A2(n4801), .A3(n4800), .A4(n4799), .ZN(n4803) );
  AOI21D0 U135 ( .A1(n4955), .A2(n4954), .B(n6856), .ZN(n4956) );
  ND4D0 U136 ( .A1(n6503), .A2(n6502), .A3(n6501), .A4(n6500), .ZN(n6509) );
  ND4D0 U137 ( .A1(n6421), .A2(n6420), .A3(n6419), .A4(n6418), .ZN(n6422) );
  ND4D0 U138 ( .A1(n6657), .A2(n6656), .A3(n6655), .A4(n6654), .ZN(n6670) );
  ND4D0 U139 ( .A1(n6575), .A2(n6574), .A3(n6573), .A4(n6572), .ZN(n6581) );
  AOI22D0 U140 ( .A1(n6914), .A2(\mem[197][1] ), .B1(n6982), .B2(\mem[194][1] ), .ZN(n6920) );
  AOI22D0 U141 ( .A1(n6872), .A2(\mem[198][1] ), .B1(n6871), .B2(\mem[249][1] ), .ZN(n6876) );
  AOI22D0 U142 ( .A1(n6914), .A2(\mem[5][1] ), .B1(n6837), .B2(\mem[15][1] ), 
        .ZN(n6838) );
  AOI22D0 U143 ( .A1(n6967), .A2(\mem[39][1] ), .B1(n6922), .B2(\mem[29][1] ), 
        .ZN(n6818) );
  AOI22D0 U144 ( .A1(n6993), .A2(\mem[181][1] ), .B1(n6916), .B2(\mem[149][1] ), .ZN(n6787) );
  AOI22D0 U145 ( .A1(n6874), .A2(\mem[170][1] ), .B1(n6995), .B2(\mem[151][1] ), .ZN(n6762) );
  ND4D0 U146 ( .A1(n5314), .A2(n5313), .A3(n5312), .A4(n5311), .ZN(n5320) );
  AOI21D0 U147 ( .A1(n6118), .A2(n6117), .B(n6856), .ZN(n6162) );
  ND4D0 U148 ( .A1(n5677), .A2(n5676), .A3(n5675), .A4(n5674), .ZN(n5688) );
  ND4D0 U149 ( .A1(n5658), .A2(n5657), .A3(n5656), .A4(n5655), .ZN(n5664) );
  AOI21D0 U150 ( .A1(n6295), .A2(n6294), .B(n6856), .ZN(n6341) );
  AOI22D0 U151 ( .A1(n6979), .A2(\mem[14][4] ), .B1(n6749), .B2(\mem[43][4] ), 
        .ZN(n185) );
  AOI22D0 U152 ( .A1(n6955), .A2(\mem[21][4] ), .B1(n6988), .B2(\mem[63][4] ), 
        .ZN(n21) );
  AOI22D0 U153 ( .A1(n6958), .A2(\mem[17][4] ), .B1(n6902), .B2(\mem[37][4] ), 
        .ZN(n5) );
  ND4D0 U154 ( .A1(n5423), .A2(n5422), .A3(n5421), .A4(n5420), .ZN(n5424) );
  ND4D0 U155 ( .A1(n5349), .A2(n5348), .A3(n5347), .A4(n5346), .ZN(n5365) );
  AOI22D0 U156 ( .A1(n6917), .A2(\mem[238][0] ), .B1(n6859), .B2(\mem[244][0] ), .ZN(n330) );
  AOI22D0 U157 ( .A1(n6979), .A2(\mem[206][0] ), .B1(n6926), .B2(\mem[193][0] ), .ZN(n317) );
  AOI22D0 U158 ( .A1(n6874), .A2(\mem[106][0] ), .B1(n6491), .B2(\mem[115][0] ), .ZN(n294) );
  AOI22D0 U159 ( .A1(n6969), .A2(\mem[82][0] ), .B1(n6869), .B2(\mem[113][0] ), 
        .ZN(n273) );
  AOI22D0 U160 ( .A1(n6861), .A2(\mem[132][0] ), .B1(n6927), .B2(\mem[153][0] ), .ZN(n250) );
  AOI22D0 U161 ( .A1(n6993), .A2(\mem[181][0] ), .B1(n6994), .B2(\mem[190][0] ), .ZN(n241) );
  AOI22D0 U162 ( .A1(n6802), .A2(\mem[152][0] ), .B1(n6979), .B2(\mem[142][0] ), .ZN(n220) );
  ND4D0 U163 ( .A1(n385), .A2(n384), .A3(n383), .A4(n382), .ZN(n386) );
  AOI22D0 U164 ( .A1(n6525), .A2(\mem[35][2] ), .B1(n6903), .B2(\mem[51][2] ), 
        .ZN(n6529) );
  AOI22D0 U165 ( .A1(n6993), .A2(\mem[53][2] ), .B1(n6994), .B2(\mem[62][2] ), 
        .ZN(n6378) );
  AOI22D0 U166 ( .A1(n6970), .A2(\mem[16][2] ), .B1(n6914), .B2(\mem[5][2] ), 
        .ZN(n6369) );
  AOI22D0 U167 ( .A1(n6892), .A2(\mem[108][3] ), .B1(n6889), .B2(\mem[92][3] ), 
        .ZN(n6701) );
  AOI22D0 U168 ( .A1(n6952), .A2(\mem[86][3] ), .B1(n6922), .B2(\mem[93][3] ), 
        .ZN(n6554) );
  ND4D0 U169 ( .A1(n6841), .A2(n6840), .A3(n6839), .A4(n6838), .ZN(n6854) );
  INVD0 U170 ( .I(n6951), .ZN(n6188) );
  ND4D0 U171 ( .A1(n182), .A2(n181), .A3(n180), .A4(n179), .ZN(n193) );
  AOI22D0 U172 ( .A1(n6639), .A2(\mem[39][5] ), .B1(n6882), .B2(\mem[15][5] ), 
        .ZN(n5485) );
  AOI22D0 U173 ( .A1(n6733), .A2(\mem[58][5] ), .B1(n6836), .B2(\mem[10][5] ), 
        .ZN(n5338) );
  AOI22D0 U174 ( .A1(n6991), .A2(\mem[20][5] ), .B1(n6174), .B2(\mem[54][5] ), 
        .ZN(n5328) );
  ND4D0 U175 ( .A1(n283), .A2(n282), .A3(n281), .A4(n280), .ZN(n299) );
  INVD0 U176 ( .I(prog_addr[1]), .ZN(n7020) );
  ND4D0 U177 ( .A1(n6529), .A2(n6528), .A3(n6527), .A4(n6526), .ZN(n6536) );
  AOI21D0 U178 ( .A1(n6649), .A2(n6648), .B(n6856), .ZN(n6696) );
  AOI22D0 U179 ( .A1(n6969), .A2(\mem[82][1] ), .B1(n6968), .B2(\mem[105][1] ), 
        .ZN(n6973) );
  AOI22D0 U180 ( .A1(n6860), .A2(\mem[99][1] ), .B1(n6774), .B2(\mem[113][1] ), 
        .ZN(n6741) );
  AOI21D0 U181 ( .A1(n5429), .A2(n5428), .B(n7004), .ZN(n5473) );
  AOI22D0 U182 ( .A1(n6914), .A2(\mem[5][0] ), .B1(n6902), .B2(\mem[37][0] ), 
        .ZN(n352) );
  AOI22D0 U183 ( .A1(n6969), .A2(\mem[18][0] ), .B1(n6874), .B2(\mem[42][0] ), 
        .ZN(n211) );
  NR2D0 U184 ( .A1(prog_addr[6]), .A2(n7527), .ZN(n7391) );
  NR2D0 U185 ( .A1(prog_addr[6]), .A2(n7458), .ZN(n7324) );
  ND4D0 U186 ( .A1(n6987), .A2(n6986), .A3(n6985), .A4(n6984), .ZN(n7001) );
  AOI211D0 U187 ( .A1(n6951), .A2(n5474), .B(n5473), .C(n5472), .ZN(n5496) );
  CKND2D0 U188 ( .A1(n7255), .A2(n7120), .ZN(n7151) );
  CKND2D0 U189 ( .A1(n7025), .A2(n7037), .ZN(n7537) );
  AOI32D0 U190 ( .A1(n6722), .A2(n6721), .A3(n6720), .B1(n7004), .B2(n6721), 
        .ZN(dout[3]) );
  INVD0 U191 ( .I(n7556), .ZN(n7557) );
  NR2D0 U192 ( .A1(n7531), .A2(n7573), .ZN(n7532) );
  INVD0 U193 ( .I(n7513), .ZN(n7514) );
  NR2D0 U194 ( .A1(n7534), .A2(n7523), .ZN(n7497) );
  INVD0 U195 ( .I(n7481), .ZN(n7482) );
  NR2D0 U196 ( .A1(n7537), .A2(n7489), .ZN(n7465) );
  INVD0 U197 ( .I(n7449), .ZN(n7450) );
  NR2D0 U198 ( .A1(n7540), .A2(n7455), .ZN(n7433) );
  INVD0 U199 ( .I(n7418), .ZN(n7419) );
  NR2D0 U200 ( .A1(n7543), .A2(n7422), .ZN(n7402) );
  INVD0 U201 ( .I(n7386), .ZN(n7387) );
  NR2D0 U202 ( .A1(n7546), .A2(n7388), .ZN(n7370) );
  INVD0 U203 ( .I(n7356), .ZN(n7357) );
  NR2D0 U204 ( .A1(n7549), .A2(n7355), .ZN(n7339) );
  INVD0 U205 ( .I(n7325), .ZN(n7326) );
  NR2D0 U206 ( .A1(n7552), .A2(n7319), .ZN(n7305) );
  INVD0 U207 ( .I(n7291), .ZN(n7292) );
  NR2D0 U208 ( .A1(n7555), .A2(n7286), .ZN(n7274) );
  INVD0 U209 ( .I(n7260), .ZN(n7261) );
  NR2D0 U210 ( .A1(n7558), .A2(n7252), .ZN(n7242) );
  INVD0 U211 ( .I(n7228), .ZN(n7229) );
  NR2D0 U212 ( .A1(n7561), .A2(n7218), .ZN(n7210) );
  INVD0 U213 ( .I(n7196), .ZN(n7197) );
  NR2D0 U214 ( .A1(n7564), .A2(n7184), .ZN(n7178) );
  INVD0 U215 ( .I(n7164), .ZN(n7165) );
  NR2D0 U216 ( .A1(n7567), .A2(n7151), .ZN(n7147) );
  INVD0 U217 ( .I(n7133), .ZN(n7134) );
  NR2D0 U218 ( .A1(n7570), .A2(n7117), .ZN(n7115) );
  INVD0 U219 ( .I(n7101), .ZN(n7102) );
  NR2D0 U220 ( .A1(n7574), .A2(n7084), .ZN(n7085) );
  INVD0 U221 ( .I(n7070), .ZN(n7071) );
  NR2D0 U222 ( .A1(n7528), .A2(n7084), .ZN(n7054) );
  INVD0 U223 ( .I(n7033), .ZN(n7034) );
  NR2D0 U224 ( .A1(n7050), .A2(n7531), .ZN(n7010) );
  NR2D0 U225 ( .A1(n7528), .A2(n7050), .ZN(n7008) );
  INVD0 U226 ( .I(addr[5]), .ZN(n13) );
  ND3D0 U227 ( .A1(addr[3]), .A2(addr[4]), .A3(n13), .ZN(n53) );
  NR2D0 U228 ( .A1(addr[2]), .A2(addr[1]), .ZN(n2) );
  CKND2D0 U229 ( .A1(addr[0]), .A2(n2), .ZN(n58) );
  NR2XD0 U230 ( .A1(n53), .A2(n58), .ZN(n6847) );
  BUFFD0 U231 ( .I(n6847), .Z(n6927) );
  INVD0 U232 ( .I(addr[0]), .ZN(n15) );
  ND3D0 U233 ( .A1(addr[2]), .A2(addr[1]), .A3(n15), .ZN(n76) );
  ND3D0 U234 ( .A1(addr[5]), .A2(addr[3]), .A3(addr[4]), .ZN(n69) );
  NR2D0 U235 ( .A1(n76), .A2(n69), .ZN(n6789) );
  BUFFD0 U236 ( .I(n6789), .Z(n6994) );
  AOI22D0 U237 ( .A1(n6927), .A2(\mem[25][4] ), .B1(n6994), .B2(\mem[62][4] ), 
        .ZN(n6) );
  INR2D0 U238 ( .A1(addr[4]), .B1(addr[3]), .ZN(n8) );
  CKND2D0 U239 ( .A1(n8), .A2(n13), .ZN(n74) );
  NR2D0 U240 ( .A1(n74), .A2(n58), .ZN(n6936) );
  BUFFD0 U241 ( .I(n6936), .Z(n6958) );
  NR2D0 U242 ( .A1(addr[3]), .A2(addr[4]), .ZN(n1) );
  CKND2D0 U243 ( .A1(addr[5]), .A2(n1), .ZN(n62) );
  INR2D0 U244 ( .A1(addr[2]), .B1(addr[1]), .ZN(n16) );
  CKND2D0 U245 ( .A1(addr[0]), .A2(n16), .ZN(n64) );
  NR2D0 U246 ( .A1(n62), .A2(n64), .ZN(n6902) );
  ND3D0 U247 ( .A1(addr[0]), .A2(addr[2]), .A3(addr[1]), .ZN(n71) );
  INR2D0 U248 ( .A1(addr[3]), .B1(addr[4]), .ZN(n14) );
  CKND2D0 U249 ( .A1(addr[5]), .A2(n14), .ZN(n59) );
  NR2XD0 U250 ( .A1(n71), .A2(n59), .ZN(n6953) );
  BUFFD0 U251 ( .I(n6953), .Z(n6179) );
  CKND2D0 U252 ( .A1(n1), .A2(n13), .ZN(n70) );
  INR2D0 U253 ( .A1(addr[1]), .B1(addr[2]), .ZN(n7) );
  CKND2D0 U254 ( .A1(n7), .A2(n15), .ZN(n73) );
  NR2D0 U255 ( .A1(n70), .A2(n73), .ZN(n6698) );
  BUFFD0 U256 ( .I(n6698), .Z(n6982) );
  AOI22D0 U257 ( .A1(n6179), .A2(\mem[47][4] ), .B1(n6982), .B2(\mem[2][4] ), 
        .ZN(n4) );
  NR2D0 U258 ( .A1(n70), .A2(n58), .ZN(n6926) );
  CKND2D0 U259 ( .A1(n2), .A2(n15), .ZN(n61) );
  NR2D0 U260 ( .A1(n61), .A2(n74), .ZN(n6881) );
  AOI22D0 U261 ( .A1(n6926), .A2(\mem[1][4] ), .B1(n6881), .B2(\mem[16][4] ), 
        .ZN(n3) );
  ND4D0 U262 ( .A1(n6), .A2(n5), .A3(n4), .A4(n3), .ZN(n28) );
  CKND2D0 U263 ( .A1(addr[0]), .A2(n7), .ZN(n60) );
  NR2XD0 U264 ( .A1(n69), .A2(n60), .ZN(n6905) );
  BUFFD0 U265 ( .I(n6905), .Z(n6530) );
  NR2D0 U266 ( .A1(n53), .A2(n73), .ZN(n6842) );
  BUFFD0 U267 ( .I(n6842), .Z(n6891) );
  AOI22D0 U268 ( .A1(n6530), .A2(\mem[59][4] ), .B1(n6891), .B2(\mem[26][4] ), 
        .ZN(n12) );
  NR2XD0 U269 ( .A1(n62), .A2(n60), .ZN(n6860) );
  CKND2D0 U270 ( .A1(addr[5]), .A2(n8), .ZN(n63) );
  NR2XD0 U271 ( .A1(n76), .A2(n63), .ZN(n6992) );
  BUFFD0 U272 ( .I(n6992), .Z(n6174) );
  AOI22D0 U273 ( .A1(n6860), .A2(\mem[35][4] ), .B1(n6174), .B2(\mem[54][4] ), 
        .ZN(n11) );
  NR2XD0 U274 ( .A1(n70), .A2(n60), .ZN(n6959) );
  BUFFD0 U275 ( .I(n6959), .Z(n6907) );
  NR2XD0 U276 ( .A1(n76), .A2(n74), .ZN(n6952) );
  BUFFD0 U277 ( .I(n6952), .Z(n6614) );
  AOI22D0 U278 ( .A1(n6907), .A2(\mem[3][4] ), .B1(n6614), .B2(\mem[22][4] ), 
        .ZN(n10) );
  NR2D0 U279 ( .A1(n71), .A2(n62), .ZN(n6639) );
  BUFFD0 U280 ( .I(n6639), .Z(n6967) );
  NR2D0 U281 ( .A1(n70), .A2(n64), .ZN(n6754) );
  AOI22D0 U282 ( .A1(n6967), .A2(\mem[39][4] ), .B1(n6754), .B2(\mem[5][4] ), 
        .ZN(n9) );
  ND4D0 U283 ( .A1(n12), .A2(n11), .A3(n10), .A4(n9), .ZN(n27) );
  NR2D0 U284 ( .A1(n61), .A2(n63), .ZN(n6983) );
  BUFFD0 U285 ( .I(n6983), .Z(n6883) );
  NR2D0 U286 ( .A1(n61), .A2(n69), .ZN(n6912) );
  AOI22D0 U287 ( .A1(n6883), .A2(\mem[48][4] ), .B1(n6912), .B2(\mem[56][4] ), 
        .ZN(n20) );
  CKND2D0 U288 ( .A1(n14), .A2(n13), .ZN(n75) );
  NR2D0 U289 ( .A1(n61), .A2(n75), .ZN(n6563) );
  NR2D0 U290 ( .A1(n71), .A2(n75), .ZN(n6837) );
  AOI22D0 U291 ( .A1(n6563), .A2(\mem[8][4] ), .B1(n6837), .B2(\mem[15][4] ), 
        .ZN(n19) );
  CKND2D0 U292 ( .A1(n16), .A2(n15), .ZN(n72) );
  NR2D0 U293 ( .A1(n72), .A2(n70), .ZN(n6835) );
  BUFFD0 U294 ( .I(n6835), .Z(n6861) );
  NR2D0 U295 ( .A1(n76), .A2(n53), .ZN(n6873) );
  BUFFD0 U296 ( .I(n6873), .Z(n6964) );
  AOI22D0 U297 ( .A1(n6861), .A2(\mem[4][4] ), .B1(n6964), .B2(\mem[30][4] ), 
        .ZN(n18) );
  NR2XD0 U298 ( .A1(n69), .A2(n64), .ZN(n6980) );
  NR2XD0 U299 ( .A1(n62), .A2(n58), .ZN(n6933) );
  AOI22D0 U300 ( .A1(n6980), .A2(\mem[61][4] ), .B1(n6933), .B2(\mem[33][4] ), 
        .ZN(n17) );
  ND4D0 U301 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NR2XD0 U302 ( .A1(n75), .A2(n58), .ZN(n6901) );
  BUFFD0 U303 ( .I(n6901), .Z(n6809) );
  NR2XD0 U304 ( .A1(n59), .A2(n73), .ZN(n6874) );
  AOI22D0 U305 ( .A1(n6809), .A2(\mem[9][4] ), .B1(n6874), .B2(\mem[42][4] ), 
        .ZN(n24) );
  NR2D0 U306 ( .A1(n72), .A2(n69), .ZN(n6870) );
  BUFFD0 U307 ( .I(n6870), .Z(n6981) );
  BUFFD0 U308 ( .I(n5966), .Z(n6680) );
  AOI22D0 U309 ( .A1(n6981), .A2(\mem[60][4] ), .B1(n6680), .B2(\mem[31][4] ), 
        .ZN(n23) );
  NR2XD0 U310 ( .A1(n72), .A2(n63), .ZN(n6728) );
  NR2D0 U311 ( .A1(n60), .A2(n74), .ZN(n6804) );
  AOI22D0 U312 ( .A1(n6728), .A2(\mem[52][4] ), .B1(n6804), .B2(\mem[19][4] ), 
        .ZN(n22) );
  NR2D0 U313 ( .A1(n64), .A2(n74), .ZN(n6916) );
  BUFFD0 U314 ( .I(n6916), .Z(n6955) );
  NR2D0 U315 ( .A1(n71), .A2(n69), .ZN(n6935) );
  BUFFD0 U316 ( .I(n6935), .Z(n6988) );
  ND4D0 U317 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NR4D0 U318 ( .A1(n28), .A2(n27), .A3(n26), .A4(n25), .ZN(n197) );
  INVD0 U319 ( .I(addr[7]), .ZN(n127) );
  NR2D0 U320 ( .A1(n127), .A2(addr[6]), .ZN(n6951) );
  NR2XD0 U321 ( .A1(n76), .A2(n70), .ZN(n6989) );
  NR2D0 U322 ( .A1(n72), .A2(n75), .ZN(n6990) );
  AOI22D0 U323 ( .A1(n6989), .A2(\mem[134][4] ), .B1(n6990), .B2(\mem[140][4] ), .ZN(n32) );
  AOI22D0 U324 ( .A1(n6983), .A2(\mem[176][4] ), .B1(n6680), .B2(\mem[159][4] ), .ZN(n31) );
  BUFFD0 U325 ( .I(n6837), .Z(n6882) );
  AOI22D0 U326 ( .A1(n6994), .A2(\mem[190][4] ), .B1(n6882), .B2(\mem[143][4] ), .ZN(n30) );
  BUFFD0 U327 ( .I(n6902), .Z(n6738) );
  AOI22D0 U328 ( .A1(n6804), .A2(\mem[147][4] ), .B1(n6738), .B2(\mem[165][4] ), .ZN(n29) );
  ND4D0 U329 ( .A1(n32), .A2(n31), .A3(n30), .A4(n29), .ZN(n48) );
  NR2XD0 U330 ( .A1(n53), .A2(n64), .ZN(n6922) );
  NR2D0 U331 ( .A1(n59), .A2(n61), .ZN(n6862) );
  AOI22D0 U332 ( .A1(n6922), .A2(\mem[157][4] ), .B1(n6862), .B2(\mem[168][4] ), .ZN(n36) );
  NR2XD0 U333 ( .A1(n59), .A2(n60), .ZN(n6868) );
  BUFFD0 U334 ( .I(n6868), .Z(n6749) );
  NR2D0 U335 ( .A1(n69), .A2(n58), .ZN(n6871) );
  BUFFD0 U336 ( .I(n6871), .Z(n6957) );
  AOI22D0 U337 ( .A1(n6749), .A2(\mem[171][4] ), .B1(n6957), .B2(\mem[185][4] ), .ZN(n35) );
  NR2D0 U338 ( .A1(n62), .A2(n76), .ZN(n6829) );
  BUFFD0 U339 ( .I(n6829), .Z(n6971) );
  NR2D0 U340 ( .A1(n63), .A2(n73), .ZN(n6966) );
  BUFFD0 U341 ( .I(n6966), .Z(n6658) );
  AOI22D0 U342 ( .A1(n6971), .A2(\mem[166][4] ), .B1(n6658), .B2(\mem[178][4] ), .ZN(n34) );
  BUFFD0 U343 ( .I(n6728), .Z(n6859) );
  AOI22D0 U344 ( .A1(n6859), .A2(\mem[180][4] ), .B1(n6174), .B2(\mem[182][4] ), .ZN(n33) );
  ND4D0 U345 ( .A1(n36), .A2(n35), .A3(n34), .A4(n33), .ZN(n47) );
  NR2XD0 U346 ( .A1(n71), .A2(n63), .ZN(n6863) );
  BUFFD0 U347 ( .I(n6863), .Z(n6803) );
  NR2D0 U348 ( .A1(n64), .A2(n75), .ZN(n6915) );
  AOI22D0 U349 ( .A1(n6803), .A2(\mem[183][4] ), .B1(n6915), .B2(\mem[141][4] ), .ZN(n40) );
  NR2D0 U350 ( .A1(n75), .A2(n73), .ZN(n6836) );
  AOI22D0 U351 ( .A1(n6980), .A2(\mem[189][4] ), .B1(n6836), .B2(\mem[138][4] ), .ZN(n39) );
  BUFFD0 U352 ( .I(n6926), .Z(n6814) );
  NR2XD0 U353 ( .A1(n62), .A2(n73), .ZN(n6923) );
  AOI22D0 U354 ( .A1(n6814), .A2(\mem[129][4] ), .B1(n6923), .B2(\mem[162][4] ), .ZN(n38) );
  AOI22D0 U355 ( .A1(n6958), .A2(\mem[145][4] ), .B1(n6563), .B2(\mem[136][4] ), .ZN(n37) );
  ND4D0 U356 ( .A1(n40), .A2(n39), .A3(n38), .A4(n37), .ZN(n46) );
  NR2XD0 U357 ( .A1(n62), .A2(n72), .ZN(n6890) );
  AOI22D0 U358 ( .A1(n6890), .A2(\mem[164][4] ), .B1(n6981), .B2(\mem[188][4] ), .ZN(n44) );
  NR2XD0 U359 ( .A1(n61), .A2(n70), .ZN(n6888) );
  NR2D0 U360 ( .A1(n58), .A2(n63), .ZN(n6869) );
  BUFFD0 U361 ( .I(n6869), .Z(n6774) );
  NR2XD0 U362 ( .A1(n59), .A2(n76), .ZN(n6917) );
  BUFFD0 U363 ( .I(n6917), .Z(n6165) );
  NR2D0 U364 ( .A1(n72), .A2(n53), .ZN(n6889) );
  AOI22D0 U365 ( .A1(n6165), .A2(\mem[174][4] ), .B1(n6889), .B2(\mem[156][4] ), .ZN(n42) );
  NR2D0 U366 ( .A1(n60), .A2(n63), .ZN(n6491) );
  AOI22D0 U367 ( .A1(n6861), .A2(\mem[132][4] ), .B1(n6491), .B2(\mem[179][4] ), .ZN(n41) );
  ND4D0 U368 ( .A1(n44), .A2(n43), .A3(n42), .A4(n41), .ZN(n45) );
  NR4D0 U369 ( .A1(n48), .A2(n47), .A3(n46), .A4(n45), .ZN(n86) );
  NR2XD0 U370 ( .A1(n53), .A2(n60), .ZN(n6913) );
  BUFFD0 U371 ( .I(n6913), .Z(n6790) );
  AOI22D0 U372 ( .A1(n6790), .A2(\mem[155][4] ), .B1(n6982), .B2(\mem[130][4] ), .ZN(n52) );
  BUFFD0 U373 ( .I(n6754), .Z(n6914) );
  AOI22D0 U374 ( .A1(n6967), .A2(\mem[167][4] ), .B1(n6914), .B2(\mem[133][4] ), .ZN(n51) );
  AOI22D0 U375 ( .A1(n6874), .A2(\mem[170][4] ), .B1(n6873), .B2(\mem[158][4] ), .ZN(n50) );
  NR2D0 U376 ( .A1(n59), .A2(n64), .ZN(n6925) );
  BUFFD0 U377 ( .I(n6925), .Z(n6760) );
  AOI22D0 U378 ( .A1(n6927), .A2(\mem[153][4] ), .B1(n6760), .B2(\mem[173][4] ), .ZN(n49) );
  ND4D0 U379 ( .A1(n52), .A2(n51), .A3(n50), .A4(n49), .ZN(n84) );
  NR2XD0 U380 ( .A1(n59), .A2(n72), .ZN(n6892) );
  NR2D0 U381 ( .A1(n71), .A2(n74), .ZN(n6707) );
  BUFFD0 U382 ( .I(n6707), .Z(n6995) );
  AOI22D0 U383 ( .A1(n6892), .A2(\mem[172][4] ), .B1(n6995), .B2(\mem[151][4] ), .ZN(n57) );
  NR2D0 U384 ( .A1(n61), .A2(n53), .ZN(n6934) );
  BUFFD0 U385 ( .I(n6934), .Z(n6802) );
  AOI22D0 U386 ( .A1(n6802), .A2(\mem[152][4] ), .B1(n6905), .B2(\mem[187][4] ), .ZN(n56) );
  BUFFD0 U387 ( .I(n6860), .Z(n6525) );
  AOI22D0 U388 ( .A1(n6525), .A2(\mem[163][4] ), .B1(n6988), .B2(\mem[191][4] ), .ZN(n55) );
  AOI22D0 U389 ( .A1(n6959), .A2(\mem[131][4] ), .B1(n6955), .B2(\mem[149][4] ), .ZN(n54) );
  ND4D0 U390 ( .A1(n57), .A2(n56), .A3(n55), .A4(n54), .ZN(n83) );
  NR2D0 U391 ( .A1(n59), .A2(n58), .ZN(n6748) );
  AOI22D0 U392 ( .A1(n6748), .A2(\mem[169][4] ), .B1(n6912), .B2(\mem[184][4] ), .ZN(n68) );
  NR2XD0 U393 ( .A1(n60), .A2(n75), .ZN(n6880) );
  AOI22D0 U394 ( .A1(n6179), .A2(\mem[175][4] ), .B1(n6880), .B2(\mem[139][4] ), .ZN(n67) );
  NR2D0 U395 ( .A1(n62), .A2(n61), .ZN(n6791) );
  BUFFD0 U396 ( .I(n6791), .Z(n6924) );
  AOI22D0 U397 ( .A1(n6901), .A2(\mem[137][4] ), .B1(n6924), .B2(\mem[160][4] ), .ZN(n66) );
  BUFFD0 U398 ( .I(n6933), .Z(n6977) );
  NR2XD0 U399 ( .A1(n64), .A2(n63), .ZN(n6993) );
  BUFFD0 U400 ( .I(n6993), .Z(n6659) );
  AOI22D0 U401 ( .A1(n6977), .A2(\mem[161][4] ), .B1(n6659), .B2(\mem[181][4] ), .ZN(n65) );
  ND4D0 U402 ( .A1(n68), .A2(n67), .A3(n66), .A4(n65), .ZN(n82) );
  BUFFD0 U403 ( .I(n6881), .Z(n6970) );
  NR2D0 U404 ( .A1(n69), .A2(n73), .ZN(n6733) );
  BUFFD0 U405 ( .I(n6733), .Z(n6879) );
  NR2XD0 U406 ( .A1(n71), .A2(n70), .ZN(n6928) );
  AOI22D0 U407 ( .A1(n6928), .A2(\mem[135][4] ), .B1(n6842), .B2(\mem[154][4] ), .ZN(n79) );
  NR2XD0 U408 ( .A1(n72), .A2(n74), .ZN(n6991) );
  NR2D0 U409 ( .A1(n74), .A2(n73), .ZN(n6542) );
  AOI22D0 U410 ( .A1(n6991), .A2(\mem[148][4] ), .B1(n6542), .B2(\mem[146][4] ), .ZN(n78) );
  NR2XD0 U411 ( .A1(n76), .A2(n75), .ZN(n6979) );
  AOI22D0 U412 ( .A1(n6979), .A2(\mem[142][4] ), .B1(n6952), .B2(\mem[150][4] ), .ZN(n77) );
  ND4D0 U413 ( .A1(n80), .A2(n79), .A3(n78), .A4(n77), .ZN(n81) );
  NR4D0 U414 ( .A1(n84), .A2(n83), .A3(n82), .A4(n81), .ZN(n85) );
  CKND2D0 U415 ( .A1(n86), .A2(n85), .ZN(n174) );
  AOI22D0 U416 ( .A1(n6989), .A2(\mem[70][4] ), .B1(n6964), .B2(\mem[94][4] ), 
        .ZN(n90) );
  AOI22D0 U417 ( .A1(n6979), .A2(\mem[78][4] ), .B1(n6680), .B2(\mem[95][4] ), 
        .ZN(n89) );
  AOI22D0 U418 ( .A1(n6861), .A2(\mem[68][4] ), .B1(n6874), .B2(\mem[106][4] ), 
        .ZN(n88) );
  AOI22D0 U419 ( .A1(n6802), .A2(\mem[88][4] ), .B1(n6791), .B2(\mem[96][4] ), 
        .ZN(n87) );
  ND4D0 U420 ( .A1(n90), .A2(n89), .A3(n88), .A4(n87), .ZN(n106) );
  AOI22D0 U421 ( .A1(n6981), .A2(\mem[124][4] ), .B1(n6888), .B2(\mem[64][4] ), 
        .ZN(n94) );
  BUFFD0 U422 ( .I(n6892), .Z(n6775) );
  AOI22D0 U423 ( .A1(n6775), .A2(\mem[108][4] ), .B1(n6912), .B2(\mem[120][4] ), .ZN(n93) );
  AOI22D0 U424 ( .A1(n6928), .A2(\mem[71][4] ), .B1(n6804), .B2(\mem[83][4] ), 
        .ZN(n92) );
  BUFFD0 U425 ( .I(n6491), .Z(n6903) );
  AOI22D0 U426 ( .A1(n6903), .A2(\mem[115][4] ), .B1(n6958), .B2(\mem[81][4] ), 
        .ZN(n91) );
  ND4D0 U427 ( .A1(n94), .A2(n93), .A3(n92), .A4(n91), .ZN(n105) );
  BUFFD0 U428 ( .I(n6990), .Z(n6906) );
  AOI22D0 U429 ( .A1(n6179), .A2(\mem[111][4] ), .B1(n6906), .B2(\mem[76][4] ), 
        .ZN(n98) );
  BUFFD0 U430 ( .I(n6889), .Z(n6784) );
  AOI22D0 U431 ( .A1(n6784), .A2(\mem[92][4] ), .B1(n6914), .B2(\mem[69][4] ), 
        .ZN(n97) );
  AOI22D0 U432 ( .A1(n6891), .A2(\mem[90][4] ), .B1(n6659), .B2(\mem[117][4] ), 
        .ZN(n96) );
  ND4D0 U433 ( .A1(n98), .A2(n97), .A3(n96), .A4(n95), .ZN(n104) );
  AOI22D0 U434 ( .A1(n6860), .A2(\mem[99][4] ), .B1(n6847), .B2(\mem[89][4] ), 
        .ZN(n102) );
  AOI22D0 U435 ( .A1(n6970), .A2(\mem[80][4] ), .B1(n6863), .B2(\mem[119][4] ), 
        .ZN(n101) );
  BUFFD0 U436 ( .I(n6991), .Z(n6747) );
  AOI22D0 U437 ( .A1(n6747), .A2(\mem[84][4] ), .B1(n6994), .B2(\mem[126][4] ), 
        .ZN(n100) );
  AOI22D0 U438 ( .A1(n6728), .A2(\mem[116][4] ), .B1(n6174), .B2(\mem[118][4] ), .ZN(n99) );
  ND4D0 U439 ( .A1(n102), .A2(n101), .A3(n100), .A4(n99), .ZN(n103) );
  NR4D0 U440 ( .A1(n106), .A2(n105), .A3(n104), .A4(n103), .ZN(n129) );
  AOI22D0 U441 ( .A1(n6809), .A2(\mem[73][4] ), .B1(n6871), .B2(\mem[121][4] ), 
        .ZN(n110) );
  BUFFD0 U442 ( .I(n6748), .Z(n6968) );
  AOI22D0 U443 ( .A1(n6968), .A2(\mem[105][4] ), .B1(n6925), .B2(\mem[109][4] ), .ZN(n109) );
  AOI22D0 U444 ( .A1(n6983), .A2(\mem[112][4] ), .B1(n6913), .B2(\mem[91][4] ), 
        .ZN(n108) );
  AOI22D0 U445 ( .A1(n6165), .A2(\mem[110][4] ), .B1(n6980), .B2(\mem[125][4] ), .ZN(n107) );
  ND4D0 U446 ( .A1(n110), .A2(n109), .A3(n108), .A4(n107), .ZN(n126) );
  BUFFD0 U447 ( .I(n6880), .Z(n6325) );
  AOI22D0 U448 ( .A1(n6325), .A2(\mem[75][4] ), .B1(n6915), .B2(\mem[77][4] ), 
        .ZN(n114) );
  AOI22D0 U449 ( .A1(n6933), .A2(\mem[97][4] ), .B1(n6542), .B2(\mem[82][4] ), 
        .ZN(n113) );
  BUFFD0 U450 ( .I(n6862), .Z(n6956) );
  AOI22D0 U451 ( .A1(n6955), .A2(\mem[85][4] ), .B1(n6956), .B2(\mem[104][4] ), 
        .ZN(n112) );
  BUFFD0 U452 ( .I(n6923), .Z(n6976) );
  AOI22D0 U453 ( .A1(n6976), .A2(\mem[98][4] ), .B1(n6698), .B2(\mem[66][4] ), 
        .ZN(n111) );
  ND4D0 U454 ( .A1(n114), .A2(n113), .A3(n112), .A4(n111), .ZN(n125) );
  AOI22D0 U455 ( .A1(n6614), .A2(\mem[86][4] ), .B1(n6774), .B2(\mem[113][4] ), 
        .ZN(n118) );
  BUFFD0 U456 ( .I(n6890), .Z(n6773) );
  BUFFD0 U457 ( .I(n6836), .Z(n6954) );
  AOI22D0 U458 ( .A1(n6773), .A2(\mem[100][4] ), .B1(n6954), .B2(\mem[74][4] ), 
        .ZN(n117) );
  BUFFD0 U459 ( .I(n6922), .Z(n6296) );
  AOI22D0 U460 ( .A1(n6733), .A2(\mem[122][4] ), .B1(n6296), .B2(\mem[93][4] ), 
        .ZN(n115) );
  AOI22D0 U461 ( .A1(n6749), .A2(\mem[107][4] ), .B1(n6563), .B2(\mem[72][4] ), 
        .ZN(n122) );
  AOI22D0 U462 ( .A1(n6967), .A2(\mem[103][4] ), .B1(n6966), .B2(\mem[114][4] ), .ZN(n121) );
  AOI22D0 U463 ( .A1(n6905), .A2(\mem[123][4] ), .B1(n6829), .B2(\mem[102][4] ), .ZN(n120) );
  AOI22D0 U464 ( .A1(n6814), .A2(\mem[65][4] ), .B1(n6935), .B2(\mem[127][4] ), 
        .ZN(n119) );
  ND4D0 U465 ( .A1(n122), .A2(n121), .A3(n120), .A4(n119), .ZN(n123) );
  NR4D0 U466 ( .A1(n126), .A2(n125), .A3(n124), .A4(n123), .ZN(n128) );
  CKND2D0 U467 ( .A1(n127), .A2(addr[6]), .ZN(n7004) );
  AOI21D0 U468 ( .A1(n129), .A2(n128), .B(n7004), .ZN(n173) );
  AOI22D0 U469 ( .A1(n6901), .A2(\mem[201][4] ), .B1(n6902), .B2(\mem[229][4] ), .ZN(n133) );
  AOI22D0 U470 ( .A1(n6954), .A2(\mem[202][4] ), .B1(n6988), .B2(\mem[255][4] ), .ZN(n132) );
  AOI22D0 U471 ( .A1(n6976), .A2(\mem[226][4] ), .B1(n6791), .B2(\mem[224][4] ), .ZN(n131) );
  AOI22D0 U472 ( .A1(n6733), .A2(\mem[250][4] ), .B1(n6804), .B2(\mem[211][4] ), .ZN(n130) );
  ND4D0 U473 ( .A1(n133), .A2(n132), .A3(n131), .A4(n130), .ZN(n149) );
  AOI22D0 U474 ( .A1(n6905), .A2(\mem[251][4] ), .B1(n6847), .B2(\mem[217][4] ), .ZN(n137) );
  AOI22D0 U475 ( .A1(n6614), .A2(\mem[214][4] ), .B1(n6956), .B2(\mem[232][4] ), .ZN(n136) );
  AOI22D0 U476 ( .A1(n6165), .A2(\mem[238][4] ), .B1(n6983), .B2(\mem[240][4] ), .ZN(n135) );
  AOI22D0 U477 ( .A1(n6784), .A2(\mem[220][4] ), .B1(n6296), .B2(\mem[221][4] ), .ZN(n134) );
  ND4D0 U478 ( .A1(n137), .A2(n136), .A3(n135), .A4(n134), .ZN(n148) );
  AOI22D0 U479 ( .A1(n6870), .A2(\mem[252][4] ), .B1(n6842), .B2(\mem[218][4] ), .ZN(n141) );
  BUFFD0 U480 ( .I(n6563), .Z(n6978) );
  AOI22D0 U481 ( .A1(n6993), .A2(\mem[245][4] ), .B1(n6978), .B2(\mem[200][4] ), .ZN(n139) );
  AOI22D0 U482 ( .A1(n6970), .A2(\mem[208][4] ), .B1(n6914), .B2(\mem[197][4] ), .ZN(n138) );
  ND4D0 U483 ( .A1(n141), .A2(n140), .A3(n139), .A4(n138), .ZN(n147) );
  AOI22D0 U484 ( .A1(n6749), .A2(\mem[235][4] ), .B1(n6990), .B2(\mem[204][4] ), .ZN(n145) );
  AOI22D0 U485 ( .A1(n6863), .A2(\mem[247][4] ), .B1(n6994), .B2(\mem[254][4] ), .ZN(n144) );
  AOI22D0 U486 ( .A1(n6707), .A2(\mem[215][4] ), .B1(n6958), .B2(\mem[209][4] ), .ZN(n143) );
  AOI22D0 U487 ( .A1(n6959), .A2(\mem[195][4] ), .B1(n6926), .B2(\mem[193][4] ), .ZN(n142) );
  ND4D0 U488 ( .A1(n145), .A2(n144), .A3(n143), .A4(n142), .ZN(n146) );
  NR4D0 U489 ( .A1(n149), .A2(n148), .A3(n147), .A4(n146), .ZN(n171) );
  BUFFD0 U490 ( .I(n6980), .Z(n6819) );
  AOI22D0 U491 ( .A1(n6819), .A2(\mem[253][4] ), .B1(n6933), .B2(\mem[225][4] ), .ZN(n153) );
  AOI22D0 U492 ( .A1(n6860), .A2(\mem[227][4] ), .B1(n6982), .B2(\mem[194][4] ), .ZN(n152) );
  AOI22D0 U493 ( .A1(n6890), .A2(\mem[228][4] ), .B1(n6913), .B2(\mem[219][4] ), .ZN(n151) );
  AOI22D0 U494 ( .A1(n6179), .A2(\mem[239][4] ), .B1(n6892), .B2(\mem[236][4] ), .ZN(n150) );
  ND4D0 U495 ( .A1(n153), .A2(n152), .A3(n151), .A4(n150), .ZN(n169) );
  AOI22D0 U496 ( .A1(n6928), .A2(\mem[199][4] ), .B1(n6979), .B2(\mem[206][4] ), .ZN(n157) );
  AOI22D0 U497 ( .A1(n6903), .A2(\mem[243][4] ), .B1(n6869), .B2(\mem[241][4] ), .ZN(n156) );
  AOI22D0 U498 ( .A1(n6971), .A2(\mem[230][4] ), .B1(n6542), .B2(\mem[210][4] ), .ZN(n155) );
  AOI22D0 U499 ( .A1(n6658), .A2(\mem[242][4] ), .B1(n6882), .B2(\mem[207][4] ), .ZN(n154) );
  ND4D0 U500 ( .A1(n157), .A2(n156), .A3(n155), .A4(n154), .ZN(n168) );
  BUFFD0 U501 ( .I(n6912), .Z(n6828) );
  AOI22D0 U502 ( .A1(n6861), .A2(\mem[196][4] ), .B1(n6828), .B2(\mem[248][4] ), .ZN(n160) );
  AOI22D0 U503 ( .A1(n6325), .A2(\mem[203][4] ), .B1(n6873), .B2(\mem[222][4] ), .ZN(n159) );
  AOI22D0 U504 ( .A1(n6888), .A2(\mem[192][4] ), .B1(n6955), .B2(\mem[213][4] ), .ZN(n158) );
  ND4D0 U505 ( .A1(n161), .A2(n160), .A3(n159), .A4(n158), .ZN(n167) );
  AOI22D0 U506 ( .A1(n6934), .A2(\mem[216][4] ), .B1(n6991), .B2(\mem[212][4] ), .ZN(n165) );
  AOI22D0 U507 ( .A1(n6680), .A2(\mem[223][4] ), .B1(n6174), .B2(\mem[246][4] ), .ZN(n164) );
  AOI22D0 U508 ( .A1(n6989), .A2(\mem[198][4] ), .B1(n6639), .B2(\mem[231][4] ), .ZN(n163) );
  AOI22D0 U509 ( .A1(n6874), .A2(\mem[234][4] ), .B1(n6957), .B2(\mem[249][4] ), .ZN(n162) );
  ND4D0 U510 ( .A1(n165), .A2(n164), .A3(n163), .A4(n162), .ZN(n166) );
  NR4D0 U511 ( .A1(n169), .A2(n168), .A3(n167), .A4(n166), .ZN(n170) );
  CKND2D0 U512 ( .A1(addr[6]), .A2(addr[7]), .ZN(n6945) );
  AOI21D0 U513 ( .A1(n171), .A2(n170), .B(n6945), .ZN(n172) );
  AOI211D0 U514 ( .A1(n6951), .A2(n174), .B(n173), .C(n172), .ZN(n196) );
  AOI22D0 U515 ( .A1(n6976), .A2(\mem[34][4] ), .B1(n6869), .B2(\mem[49][4] ), 
        .ZN(n178) );
  AOI22D0 U516 ( .A1(n6971), .A2(\mem[38][4] ), .B1(n6836), .B2(\mem[10][4] ), 
        .ZN(n177) );
  AOI22D0 U517 ( .A1(n6790), .A2(\mem[27][4] ), .B1(n6925), .B2(\mem[45][4] ), 
        .ZN(n176) );
  AOI22D0 U518 ( .A1(n6890), .A2(\mem[36][4] ), .B1(n6889), .B2(\mem[28][4] ), 
        .ZN(n175) );
  ND4D0 U519 ( .A1(n178), .A2(n177), .A3(n176), .A4(n175), .ZN(n194) );
  AOI22D0 U520 ( .A1(n6968), .A2(\mem[41][4] ), .B1(n6906), .B2(\mem[12][4] ), 
        .ZN(n182) );
  BUFFD0 U521 ( .I(n6989), .Z(n6872) );
  AOI22D0 U522 ( .A1(n6872), .A2(\mem[6][4] ), .B1(n6888), .B2(\mem[0][4] ), 
        .ZN(n181) );
  AOI22D0 U523 ( .A1(n6892), .A2(\mem[44][4] ), .B1(n6903), .B2(\mem[51][4] ), 
        .ZN(n180) );
  BUFFD0 U524 ( .I(n6915), .Z(n6965) );
  AOI22D0 U525 ( .A1(n6863), .A2(\mem[55][4] ), .B1(n6965), .B2(\mem[13][4] ), 
        .ZN(n179) );
  AOI22D0 U526 ( .A1(n6879), .A2(\mem[58][4] ), .B1(n6658), .B2(\mem[50][4] ), 
        .ZN(n186) );
  AOI22D0 U527 ( .A1(n6165), .A2(\mem[46][4] ), .B1(n6871), .B2(\mem[57][4] ), 
        .ZN(n184) );
  BUFFD0 U528 ( .I(n6542), .Z(n6969) );
  AOI22D0 U529 ( .A1(n6991), .A2(\mem[20][4] ), .B1(n6969), .B2(\mem[18][4] ), 
        .ZN(n183) );
  ND4D0 U530 ( .A1(n186), .A2(n185), .A3(n184), .A4(n183), .ZN(n192) );
  AOI22D0 U531 ( .A1(n6993), .A2(\mem[53][4] ), .B1(n6862), .B2(\mem[40][4] ), 
        .ZN(n190) );
  BUFFD0 U532 ( .I(n6928), .Z(n6830) );
  AOI22D0 U533 ( .A1(n6830), .A2(\mem[7][4] ), .B1(n6880), .B2(\mem[11][4] ), 
        .ZN(n189) );
  AOI22D0 U534 ( .A1(n6922), .A2(\mem[29][4] ), .B1(n6995), .B2(\mem[23][4] ), 
        .ZN(n188) );
  AOI22D0 U535 ( .A1(n6802), .A2(\mem[24][4] ), .B1(n6924), .B2(\mem[32][4] ), 
        .ZN(n187) );
  ND4D0 U536 ( .A1(n190), .A2(n189), .A3(n188), .A4(n187), .ZN(n191) );
  NR4D0 U537 ( .A1(n194), .A2(n193), .A3(n192), .A4(n191), .ZN(n195) );
  OR2D0 U538 ( .A1(addr[6]), .A2(addr[7]), .Z(n6856) );
  AOI32D0 U539 ( .A1(n197), .A2(n196), .A3(n195), .B1(n6856), .B2(n196), .ZN(
        dout[4]) );
  AOI22D0 U540 ( .A1(n6977), .A2(\mem[33][0] ), .B1(n6835), .B2(\mem[4][0] ), 
        .ZN(n201) );
  AOI22D0 U541 ( .A1(n6879), .A2(\mem[58][0] ), .B1(n6954), .B2(\mem[10][0] ), 
        .ZN(n200) );
  AOI22D0 U542 ( .A1(n6802), .A2(\mem[24][0] ), .B1(n6901), .B2(\mem[9][0] ), 
        .ZN(n199) );
  AOI22D0 U543 ( .A1(n6784), .A2(\mem[28][0] ), .B1(n6829), .B2(\mem[38][0] ), 
        .ZN(n198) );
  ND4D0 U544 ( .A1(n201), .A2(n200), .A3(n199), .A4(n198), .ZN(n217) );
  AOI22D0 U545 ( .A1(n6928), .A2(\mem[7][0] ), .B1(n6860), .B2(\mem[35][0] ), 
        .ZN(n205) );
  AOI22D0 U546 ( .A1(n6814), .A2(\mem[1][0] ), .B1(n6760), .B2(\mem[45][0] ), 
        .ZN(n204) );
  AOI22D0 U547 ( .A1(n6913), .A2(\mem[27][0] ), .B1(n6563), .B2(\mem[8][0] ), 
        .ZN(n203) );
  AOI22D0 U548 ( .A1(n6868), .A2(\mem[43][0] ), .B1(n6847), .B2(\mem[25][0] ), 
        .ZN(n202) );
  ND4D0 U549 ( .A1(n205), .A2(n204), .A3(n203), .A4(n202), .ZN(n216) );
  AOI22D0 U550 ( .A1(n6959), .A2(\mem[3][0] ), .B1(n6659), .B2(\mem[53][0] ), 
        .ZN(n209) );
  AOI22D0 U551 ( .A1(n6968), .A2(\mem[41][0] ), .B1(n6828), .B2(\mem[56][0] ), 
        .ZN(n208) );
  AOI22D0 U552 ( .A1(n6979), .A2(\mem[14][0] ), .B1(n6966), .B2(\mem[50][0] ), 
        .ZN(n207) );
  AOI22D0 U553 ( .A1(n6955), .A2(\mem[21][0] ), .B1(n6906), .B2(\mem[12][0] ), 
        .ZN(n206) );
  ND4D0 U554 ( .A1(n209), .A2(n208), .A3(n207), .A4(n206), .ZN(n215) );
  AOI22D0 U555 ( .A1(n6991), .A2(\mem[20][0] ), .B1(n6891), .B2(\mem[26][0] ), 
        .ZN(n213) );
  AOI22D0 U556 ( .A1(n6880), .A2(\mem[11][0] ), .B1(n6958), .B2(\mem[17][0] ), 
        .ZN(n212) );
  AOI22D0 U557 ( .A1(n6980), .A2(\mem[61][0] ), .B1(n6967), .B2(\mem[39][0] ), 
        .ZN(n210) );
  ND4D0 U558 ( .A1(n213), .A2(n212), .A3(n211), .A4(n210), .ZN(n214) );
  NR4D0 U559 ( .A1(n217), .A2(n216), .A3(n215), .A4(n214), .ZN(n369) );
  AOI22D0 U560 ( .A1(n6870), .A2(\mem[188][0] ), .B1(n6874), .B2(\mem[170][0] ), .ZN(n221) );
  AOI22D0 U561 ( .A1(n6814), .A2(\mem[129][0] ), .B1(n6933), .B2(\mem[161][0] ), .ZN(n219) );
  AOI22D0 U562 ( .A1(n6953), .A2(\mem[175][0] ), .B1(n6992), .B2(\mem[182][0] ), .ZN(n218) );
  ND4D0 U563 ( .A1(n221), .A2(n220), .A3(n219), .A4(n218), .ZN(n237) );
  AOI22D0 U564 ( .A1(n6989), .A2(\mem[134][0] ), .B1(n6863), .B2(\mem[183][0] ), .ZN(n225) );
  AOI22D0 U565 ( .A1(n6971), .A2(\mem[166][0] ), .B1(n6542), .B2(\mem[146][0] ), .ZN(n224) );
  AOI22D0 U566 ( .A1(n6880), .A2(\mem[139][0] ), .B1(n6774), .B2(\mem[177][0] ), .ZN(n223) );
  AOI22D0 U567 ( .A1(n6879), .A2(\mem[186][0] ), .B1(n6924), .B2(\mem[160][0] ), .ZN(n222) );
  ND4D0 U568 ( .A1(n225), .A2(n224), .A3(n223), .A4(n222), .ZN(n236) );
  AOI22D0 U569 ( .A1(n6891), .A2(\mem[154][0] ), .B1(n6871), .B2(\mem[185][0] ), .ZN(n229) );
  AOI22D0 U570 ( .A1(n6959), .A2(\mem[131][0] ), .B1(n6958), .B2(\mem[145][0] ), .ZN(n228) );
  AOI22D0 U571 ( .A1(n6773), .A2(\mem[164][0] ), .B1(n6905), .B2(\mem[187][0] ), .ZN(n227) );
  AOI22D0 U572 ( .A1(n6922), .A2(\mem[157][0] ), .B1(n6707), .B2(\mem[151][0] ), .ZN(n226) );
  ND4D0 U573 ( .A1(n229), .A2(n228), .A3(n227), .A4(n226), .ZN(n235) );
  AOI22D0 U574 ( .A1(n6968), .A2(\mem[169][0] ), .B1(n6956), .B2(\mem[168][0] ), .ZN(n233) );
  AOI22D0 U575 ( .A1(n6728), .A2(\mem[180][0] ), .B1(n6978), .B2(\mem[136][0] ), .ZN(n232) );
  AOI22D0 U576 ( .A1(n6860), .A2(\mem[163][0] ), .B1(n6738), .B2(\mem[165][0] ), .ZN(n231) );
  AOI22D0 U577 ( .A1(n6935), .A2(\mem[191][0] ), .B1(n6882), .B2(\mem[143][0] ), .ZN(n230) );
  ND4D0 U578 ( .A1(n233), .A2(n232), .A3(n231), .A4(n230), .ZN(n234) );
  NR4D0 U579 ( .A1(n237), .A2(n236), .A3(n235), .A4(n234), .ZN(n259) );
  AOI22D0 U580 ( .A1(n6614), .A2(\mem[150][0] ), .B1(n6889), .B2(\mem[156][0] ), .ZN(n240) );
  AOI22D0 U581 ( .A1(n6982), .A2(\mem[130][0] ), .B1(n6828), .B2(\mem[184][0] ), .ZN(n239) );
  AOI22D0 U582 ( .A1(n6888), .A2(\mem[128][0] ), .B1(n6790), .B2(\mem[155][0] ), .ZN(n238) );
  ND4D0 U583 ( .A1(n241), .A2(n240), .A3(n239), .A4(n238), .ZN(n257) );
  AOI22D0 U584 ( .A1(n6954), .A2(\mem[138][0] ), .B1(n6990), .B2(\mem[140][0] ), .ZN(n245) );
  AOI22D0 U585 ( .A1(n6967), .A2(\mem[167][0] ), .B1(n6914), .B2(\mem[133][0] ), .ZN(n244) );
  AOI22D0 U586 ( .A1(n6917), .A2(\mem[174][0] ), .B1(n6966), .B2(\mem[178][0] ), .ZN(n243) );
  AOI22D0 U587 ( .A1(n6970), .A2(\mem[144][0] ), .B1(n6901), .B2(\mem[137][0] ), .ZN(n242) );
  ND4D0 U588 ( .A1(n245), .A2(n244), .A3(n243), .A4(n242), .ZN(n256) );
  AOI22D0 U589 ( .A1(n6928), .A2(\mem[135][0] ), .B1(n6991), .B2(\mem[148][0] ), .ZN(n249) );
  AOI22D0 U590 ( .A1(n6892), .A2(\mem[172][0] ), .B1(n6976), .B2(\mem[162][0] ), .ZN(n248) );
  BUFFD0 U591 ( .I(n6804), .Z(n6904) );
  AOI22D0 U592 ( .A1(n6904), .A2(\mem[147][0] ), .B1(n6873), .B2(\mem[158][0] ), .ZN(n247) );
  AOI22D0 U593 ( .A1(n6749), .A2(\mem[171][0] ), .B1(n6925), .B2(\mem[173][0] ), .ZN(n246) );
  ND4D0 U594 ( .A1(n249), .A2(n248), .A3(n247), .A4(n246), .ZN(n255) );
  AOI22D0 U595 ( .A1(n6980), .A2(\mem[189][0] ), .B1(n5966), .B2(\mem[159][0] ), .ZN(n253) );
  AOI22D0 U596 ( .A1(n6903), .A2(\mem[179][0] ), .B1(n6916), .B2(\mem[149][0] ), .ZN(n252) );
  AOI22D0 U597 ( .A1(n6883), .A2(\mem[176][0] ), .B1(n6965), .B2(\mem[141][0] ), .ZN(n251) );
  ND4D0 U598 ( .A1(n253), .A2(n252), .A3(n251), .A4(n250), .ZN(n254) );
  NR4D0 U599 ( .A1(n257), .A2(n256), .A3(n255), .A4(n254), .ZN(n258) );
  CKND2D0 U600 ( .A1(n259), .A2(n258), .ZN(n346) );
  AOI22D0 U601 ( .A1(n6658), .A2(\mem[114][0] ), .B1(n6563), .B2(\mem[72][0] ), 
        .ZN(n263) );
  AOI22D0 U602 ( .A1(n6980), .A2(\mem[125][0] ), .B1(n6905), .B2(\mem[123][0] ), .ZN(n262) );
  AOI22D0 U603 ( .A1(n6917), .A2(\mem[110][0] ), .B1(n6871), .B2(\mem[121][0] ), .ZN(n261) );
  AOI22D0 U604 ( .A1(n6842), .A2(\mem[90][0] ), .B1(n6859), .B2(\mem[116][0] ), 
        .ZN(n260) );
  ND4D0 U605 ( .A1(n263), .A2(n262), .A3(n261), .A4(n260), .ZN(n279) );
  AOI22D0 U606 ( .A1(n6967), .A2(\mem[103][0] ), .B1(n6914), .B2(\mem[69][0] ), 
        .ZN(n267) );
  AOI22D0 U607 ( .A1(n6883), .A2(\mem[112][0] ), .B1(n6992), .B2(\mem[118][0] ), .ZN(n266) );
  AOI22D0 U608 ( .A1(n6958), .A2(\mem[81][0] ), .B1(n6994), .B2(\mem[126][0] ), 
        .ZN(n265) );
  AOI22D0 U609 ( .A1(n6784), .A2(\mem[92][0] ), .B1(n6935), .B2(\mem[127][0] ), 
        .ZN(n264) );
  ND4D0 U610 ( .A1(n267), .A2(n266), .A3(n265), .A4(n264), .ZN(n278) );
  AOI22D0 U611 ( .A1(n6868), .A2(\mem[107][0] ), .B1(n6888), .B2(\mem[64][0] ), 
        .ZN(n271) );
  AOI22D0 U612 ( .A1(n6861), .A2(\mem[68][0] ), .B1(n6881), .B2(\mem[80][0] ), 
        .ZN(n270) );
  AOI22D0 U613 ( .A1(n6982), .A2(\mem[66][0] ), .B1(n6956), .B2(\mem[104][0] ), 
        .ZN(n269) );
  AOI22D0 U614 ( .A1(n6928), .A2(\mem[71][0] ), .B1(n5966), .B2(\mem[95][0] ), 
        .ZN(n268) );
  ND4D0 U615 ( .A1(n271), .A2(n270), .A3(n269), .A4(n268), .ZN(n277) );
  AOI22D0 U616 ( .A1(n6890), .A2(\mem[100][0] ), .B1(n6912), .B2(\mem[120][0] ), .ZN(n275) );
  AOI22D0 U617 ( .A1(n6959), .A2(\mem[67][0] ), .B1(n6860), .B2(\mem[99][0] ), 
        .ZN(n274) );
  AOI22D0 U618 ( .A1(n6952), .A2(\mem[86][0] ), .B1(n6913), .B2(\mem[91][0] ), 
        .ZN(n272) );
  ND4D0 U619 ( .A1(n275), .A2(n274), .A3(n273), .A4(n272), .ZN(n276) );
  NR4D0 U620 ( .A1(n279), .A2(n278), .A3(n277), .A4(n276), .ZN(n301) );
  AOI22D0 U621 ( .A1(n6955), .A2(\mem[85][0] ), .B1(n6836), .B2(\mem[74][0] ), 
        .ZN(n283) );
  AOI22D0 U622 ( .A1(n6879), .A2(\mem[122][0] ), .B1(n6659), .B2(\mem[117][0] ), .ZN(n282) );
  AOI22D0 U623 ( .A1(n6979), .A2(\mem[78][0] ), .B1(n6976), .B2(\mem[98][0] ), 
        .ZN(n281) );
  AOI22D0 U624 ( .A1(n6892), .A2(\mem[108][0] ), .B1(n6837), .B2(\mem[79][0] ), 
        .ZN(n280) );
  AOI22D0 U625 ( .A1(n6847), .A2(\mem[89][0] ), .B1(n6922), .B2(\mem[93][0] ), 
        .ZN(n287) );
  AOI22D0 U626 ( .A1(n6981), .A2(\mem[124][0] ), .B1(n6738), .B2(\mem[101][0] ), .ZN(n286) );
  AOI22D0 U627 ( .A1(n6989), .A2(\mem[70][0] ), .B1(n6990), .B2(\mem[76][0] ), 
        .ZN(n285) );
  AOI22D0 U628 ( .A1(n6814), .A2(\mem[65][0] ), .B1(n6791), .B2(\mem[96][0] ), 
        .ZN(n284) );
  ND4D0 U629 ( .A1(n287), .A2(n286), .A3(n285), .A4(n284), .ZN(n298) );
  AOI22D0 U630 ( .A1(n6915), .A2(\mem[77][0] ), .B1(n6925), .B2(\mem[109][0] ), 
        .ZN(n291) );
  AOI22D0 U631 ( .A1(n6953), .A2(\mem[111][0] ), .B1(n6968), .B2(\mem[105][0] ), .ZN(n290) );
  AOI22D0 U632 ( .A1(n6991), .A2(\mem[84][0] ), .B1(n6901), .B2(\mem[73][0] ), 
        .ZN(n289) );
  AOI22D0 U633 ( .A1(n6934), .A2(\mem[88][0] ), .B1(n6977), .B2(\mem[97][0] ), 
        .ZN(n288) );
  ND4D0 U634 ( .A1(n291), .A2(n290), .A3(n289), .A4(n288), .ZN(n297) );
  AOI22D0 U635 ( .A1(n6880), .A2(\mem[75][0] ), .B1(n6829), .B2(\mem[102][0] ), 
        .ZN(n295) );
  AOI22D0 U636 ( .A1(n6995), .A2(\mem[87][0] ), .B1(n6904), .B2(\mem[83][0] ), 
        .ZN(n293) );
  AOI22D0 U637 ( .A1(n6863), .A2(\mem[119][0] ), .B1(n6873), .B2(\mem[94][0] ), 
        .ZN(n292) );
  ND4D0 U638 ( .A1(n295), .A2(n294), .A3(n293), .A4(n292), .ZN(n296) );
  NR4D0 U639 ( .A1(n299), .A2(n298), .A3(n297), .A4(n296), .ZN(n300) );
  AOI21D0 U640 ( .A1(n301), .A2(n300), .B(n7004), .ZN(n345) );
  AOI22D0 U641 ( .A1(n6967), .A2(\mem[231][0] ), .B1(n6837), .B2(\mem[207][0] ), .ZN(n305) );
  AOI22D0 U642 ( .A1(n6802), .A2(\mem[216][0] ), .B1(n6954), .B2(\mem[202][0] ), .ZN(n304) );
  AOI22D0 U643 ( .A1(n6923), .A2(\mem[226][0] ), .B1(n6925), .B2(\mem[237][0] ), .ZN(n303) );
  AOI22D0 U644 ( .A1(n6892), .A2(\mem[236][0] ), .B1(n6903), .B2(\mem[243][0] ), .ZN(n302) );
  ND4D0 U645 ( .A1(n305), .A2(n304), .A3(n303), .A4(n302), .ZN(n321) );
  AOI22D0 U646 ( .A1(n6860), .A2(\mem[227][0] ), .B1(n6881), .B2(\mem[208][0] ), .ZN(n309) );
  AOI22D0 U647 ( .A1(n6928), .A2(\mem[199][0] ), .B1(n6935), .B2(\mem[255][0] ), .ZN(n308) );
  AOI22D0 U648 ( .A1(n6862), .A2(\mem[232][0] ), .B1(n6912), .B2(\mem[248][0] ), .ZN(n307) );
  AOI22D0 U649 ( .A1(n6933), .A2(\mem[225][0] ), .B1(n6774), .B2(\mem[241][0] ), .ZN(n306) );
  ND4D0 U650 ( .A1(n309), .A2(n308), .A3(n307), .A4(n306), .ZN(n320) );
  AOI22D0 U651 ( .A1(n6905), .A2(\mem[251][0] ), .B1(n6871), .B2(\mem[249][0] ), .ZN(n313) );
  AOI22D0 U652 ( .A1(n6738), .A2(\mem[229][0] ), .B1(n6873), .B2(\mem[222][0] ), .ZN(n312) );
  AOI22D0 U653 ( .A1(n6784), .A2(\mem[220][0] ), .B1(n6891), .B2(\mem[218][0] ), .ZN(n311) );
  AOI22D0 U654 ( .A1(n6863), .A2(\mem[247][0] ), .B1(n6990), .B2(\mem[204][0] ), .ZN(n310) );
  ND4D0 U655 ( .A1(n313), .A2(n312), .A3(n311), .A4(n310), .ZN(n319) );
  AOI22D0 U656 ( .A1(n6809), .A2(\mem[201][0] ), .B1(n6915), .B2(\mem[205][0] ), .ZN(n316) );
  AOI22D0 U657 ( .A1(n6904), .A2(\mem[211][0] ), .B1(n6748), .B2(\mem[233][0] ), .ZN(n315) );
  AOI22D0 U658 ( .A1(n6861), .A2(\mem[196][0] ), .B1(n6847), .B2(\mem[217][0] ), .ZN(n314) );
  ND4D0 U659 ( .A1(n317), .A2(n316), .A3(n315), .A4(n314), .ZN(n318) );
  NR4D0 U660 ( .A1(n321), .A2(n320), .A3(n319), .A4(n318), .ZN(n343) );
  BUFFD0 U661 ( .I(n6874), .Z(n6727) );
  AOI22D0 U662 ( .A1(n6727), .A2(\mem[234][0] ), .B1(n6922), .B2(\mem[221][0] ), .ZN(n325) );
  AOI22D0 U663 ( .A1(n6880), .A2(\mem[203][0] ), .B1(n6958), .B2(\mem[209][0] ), .ZN(n324) );
  AOI22D0 U664 ( .A1(n6953), .A2(\mem[239][0] ), .B1(n6994), .B2(\mem[254][0] ), .ZN(n323) );
  AOI22D0 U665 ( .A1(n6969), .A2(\mem[210][0] ), .B1(n6680), .B2(\mem[223][0] ), .ZN(n322) );
  ND4D0 U666 ( .A1(n325), .A2(n324), .A3(n323), .A4(n322), .ZN(n341) );
  AOI22D0 U667 ( .A1(n6868), .A2(\mem[235][0] ), .B1(n6563), .B2(\mem[200][0] ), .ZN(n329) );
  AOI22D0 U668 ( .A1(n6733), .A2(\mem[250][0] ), .B1(n6955), .B2(\mem[213][0] ), .ZN(n328) );
  AOI22D0 U669 ( .A1(n6971), .A2(\mem[230][0] ), .B1(n6914), .B2(\mem[197][0] ), .ZN(n327) );
  AOI22D0 U670 ( .A1(n6959), .A2(\mem[195][0] ), .B1(n6983), .B2(\mem[240][0] ), .ZN(n326) );
  ND4D0 U671 ( .A1(n329), .A2(n328), .A3(n327), .A4(n326), .ZN(n340) );
  AOI22D0 U672 ( .A1(n6995), .A2(\mem[215][0] ), .B1(n6982), .B2(\mem[194][0] ), .ZN(n333) );
  AOI22D0 U673 ( .A1(n6890), .A2(\mem[228][0] ), .B1(n6913), .B2(\mem[219][0] ), .ZN(n332) );
  AOI22D0 U674 ( .A1(n6991), .A2(\mem[212][0] ), .B1(n6993), .B2(\mem[245][0] ), .ZN(n331) );
  ND4D0 U675 ( .A1(n333), .A2(n332), .A3(n331), .A4(n330), .ZN(n339) );
  AOI22D0 U676 ( .A1(n6989), .A2(\mem[198][0] ), .B1(n6888), .B2(\mem[192][0] ), .ZN(n337) );
  AOI22D0 U677 ( .A1(n6870), .A2(\mem[252][0] ), .B1(n6952), .B2(\mem[214][0] ), .ZN(n336) );
  AOI22D0 U678 ( .A1(n6980), .A2(\mem[253][0] ), .B1(n6924), .B2(\mem[224][0] ), .ZN(n335) );
  AOI22D0 U679 ( .A1(n6658), .A2(\mem[242][0] ), .B1(n6992), .B2(\mem[246][0] ), .ZN(n334) );
  ND4D0 U680 ( .A1(n337), .A2(n336), .A3(n335), .A4(n334), .ZN(n338) );
  NR4D0 U681 ( .A1(n341), .A2(n340), .A3(n339), .A4(n338), .ZN(n342) );
  AOI21D0 U682 ( .A1(n343), .A2(n342), .B(n6945), .ZN(n344) );
  AOI211D0 U683 ( .A1(n6951), .A2(n346), .B(n345), .C(n344), .ZN(n368) );
  AOI22D0 U684 ( .A1(n6917), .A2(\mem[46][0] ), .B1(n6923), .B2(\mem[34][0] ), 
        .ZN(n350) );
  AOI22D0 U685 ( .A1(n6892), .A2(\mem[44][0] ), .B1(n6789), .B2(\mem[62][0] ), 
        .ZN(n349) );
  AOI22D0 U686 ( .A1(n6957), .A2(\mem[57][0] ), .B1(n6992), .B2(\mem[54][0] ), 
        .ZN(n348) );
  AOI22D0 U687 ( .A1(n6863), .A2(\mem[55][0] ), .B1(n6296), .B2(\mem[29][0] ), 
        .ZN(n347) );
  ND4D0 U688 ( .A1(n350), .A2(n349), .A3(n348), .A4(n347), .ZN(n366) );
  AOI22D0 U689 ( .A1(n6791), .A2(\mem[32][0] ), .B1(n6915), .B2(\mem[13][0] ), 
        .ZN(n354) );
  AOI22D0 U690 ( .A1(n6970), .A2(\mem[16][0] ), .B1(n6888), .B2(\mem[0][0] ), 
        .ZN(n353) );
  AOI22D0 U691 ( .A1(n6952), .A2(\mem[22][0] ), .B1(n5966), .B2(\mem[31][0] ), 
        .ZN(n351) );
  ND4D0 U692 ( .A1(n354), .A2(n353), .A3(n352), .A4(n351), .ZN(n365) );
  AOI22D0 U693 ( .A1(n6905), .A2(\mem[59][0] ), .B1(n6837), .B2(\mem[15][0] ), 
        .ZN(n358) );
  AOI22D0 U694 ( .A1(n6491), .A2(\mem[51][0] ), .B1(n6935), .B2(\mem[63][0] ), 
        .ZN(n357) );
  AOI22D0 U695 ( .A1(n6870), .A2(\mem[60][0] ), .B1(n6983), .B2(\mem[48][0] ), 
        .ZN(n356) );
  AOI22D0 U696 ( .A1(n6904), .A2(\mem[19][0] ), .B1(n6869), .B2(\mem[49][0] ), 
        .ZN(n355) );
  ND4D0 U697 ( .A1(n358), .A2(n357), .A3(n356), .A4(n355), .ZN(n364) );
  AOI22D0 U698 ( .A1(n6995), .A2(\mem[23][0] ), .B1(n6698), .B2(\mem[2][0] ), 
        .ZN(n362) );
  AOI22D0 U699 ( .A1(n6989), .A2(\mem[6][0] ), .B1(n6728), .B2(\mem[52][0] ), 
        .ZN(n361) );
  AOI22D0 U700 ( .A1(n6956), .A2(\mem[40][0] ), .B1(n6873), .B2(\mem[30][0] ), 
        .ZN(n360) );
  AOI22D0 U701 ( .A1(n6953), .A2(\mem[47][0] ), .B1(n6890), .B2(\mem[36][0] ), 
        .ZN(n359) );
  ND4D0 U702 ( .A1(n362), .A2(n361), .A3(n360), .A4(n359), .ZN(n363) );
  NR4D0 U703 ( .A1(n366), .A2(n365), .A3(n364), .A4(n363), .ZN(n367) );
  AOI32D0 U704 ( .A1(n369), .A2(n368), .A3(n367), .B1(n6856), .B2(n368), .ZN(
        dout[0]) );
  AOI22D0 U705 ( .A1(n6680), .A2(\mem[95][13] ), .B1(n6491), .B2(
        \mem[115][13] ), .ZN(n373) );
  AOI22D0 U706 ( .A1(n6980), .A2(\mem[125][13] ), .B1(n6989), .B2(
        \mem[70][13] ), .ZN(n372) );
  AOI22D0 U707 ( .A1(n6883), .A2(\mem[112][13] ), .B1(n6992), .B2(
        \mem[118][13] ), .ZN(n371) );
  AOI22D0 U708 ( .A1(n6976), .A2(\mem[98][13] ), .B1(n6828), .B2(
        \mem[120][13] ), .ZN(n370) );
  ND4D0 U709 ( .A1(n373), .A2(n372), .A3(n371), .A4(n370), .ZN(n389) );
  AOI22D0 U710 ( .A1(n6934), .A2(\mem[88][13] ), .B1(n6991), .B2(\mem[84][13] ), .ZN(n377) );
  BUFFD0 U711 ( .I(n6979), .Z(n6759) );
  AOI22D0 U712 ( .A1(n6759), .A2(\mem[78][13] ), .B1(n6868), .B2(
        \mem[107][13] ), .ZN(n376) );
  AOI22D0 U713 ( .A1(n6525), .A2(\mem[99][13] ), .B1(n6774), .B2(
        \mem[113][13] ), .ZN(n375) );
  AOI22D0 U714 ( .A1(n6954), .A2(\mem[74][13] ), .B1(n6882), .B2(\mem[79][13] ), .ZN(n374) );
  ND4D0 U715 ( .A1(n377), .A2(n376), .A3(n375), .A4(n374), .ZN(n388) );
  AOI22D0 U716 ( .A1(n6890), .A2(\mem[100][13] ), .B1(n6881), .B2(
        \mem[80][13] ), .ZN(n381) );
  AOI22D0 U717 ( .A1(n6888), .A2(\mem[64][13] ), .B1(n6809), .B2(\mem[73][13] ), .ZN(n380) );
  AOI22D0 U718 ( .A1(n6969), .A2(\mem[82][13] ), .B1(n6748), .B2(
        \mem[105][13] ), .ZN(n379) );
  AOI22D0 U719 ( .A1(n6971), .A2(\mem[102][13] ), .B1(n6728), .B2(
        \mem[116][13] ), .ZN(n378) );
  ND4D0 U720 ( .A1(n381), .A2(n380), .A3(n379), .A4(n378), .ZN(n387) );
  AOI22D0 U721 ( .A1(n6727), .A2(\mem[106][13] ), .B1(n6965), .B2(
        \mem[77][13] ), .ZN(n385) );
  AOI22D0 U722 ( .A1(n6924), .A2(\mem[96][13] ), .B1(n6789), .B2(
        \mem[126][13] ), .ZN(n384) );
  AOI22D0 U723 ( .A1(n6917), .A2(\mem[110][13] ), .B1(n6964), .B2(
        \mem[94][13] ), .ZN(n382) );
  NR4D0 U724 ( .A1(n389), .A2(n388), .A3(n387), .A4(n386), .ZN(n541) );
  AOI22D0 U725 ( .A1(n6870), .A2(\mem[188][13] ), .B1(n6639), .B2(
        \mem[167][13] ), .ZN(n393) );
  AOI22D0 U726 ( .A1(n6883), .A2(\mem[176][13] ), .B1(n6738), .B2(
        \mem[165][13] ), .ZN(n392) );
  AOI22D0 U727 ( .A1(n6872), .A2(\mem[134][13] ), .B1(n6836), .B2(
        \mem[138][13] ), .ZN(n391) );
  AOI22D0 U728 ( .A1(n6980), .A2(\mem[189][13] ), .B1(n6542), .B2(
        \mem[146][13] ), .ZN(n390) );
  ND4D0 U729 ( .A1(n393), .A2(n392), .A3(n391), .A4(n390), .ZN(n409) );
  AOI22D0 U730 ( .A1(n6880), .A2(\mem[139][13] ), .B1(n6863), .B2(
        \mem[183][13] ), .ZN(n397) );
  AOI22D0 U731 ( .A1(n6922), .A2(\mem[157][13] ), .B1(n6916), .B2(
        \mem[149][13] ), .ZN(n396) );
  AOI22D0 U732 ( .A1(n6680), .A2(\mem[159][13] ), .B1(n6978), .B2(
        \mem[136][13] ), .ZN(n395) );
  AOI22D0 U733 ( .A1(n6530), .A2(\mem[187][13] ), .B1(n6882), .B2(
        \mem[143][13] ), .ZN(n394) );
  ND4D0 U734 ( .A1(n397), .A2(n396), .A3(n395), .A4(n394), .ZN(n408) );
  AOI22D0 U735 ( .A1(n6958), .A2(\mem[145][13] ), .B1(n6774), .B2(
        \mem[177][13] ), .ZN(n401) );
  AOI22D0 U736 ( .A1(n6802), .A2(\mem[152][13] ), .B1(n6698), .B2(
        \mem[130][13] ), .ZN(n400) );
  AOI22D0 U737 ( .A1(n6747), .A2(\mem[148][13] ), .B1(n6733), .B2(
        \mem[186][13] ), .ZN(n399) );
  AOI22D0 U738 ( .A1(n6933), .A2(\mem[161][13] ), .B1(n6809), .B2(
        \mem[137][13] ), .ZN(n398) );
  ND4D0 U739 ( .A1(n401), .A2(n400), .A3(n399), .A4(n398), .ZN(n407) );
  AOI22D0 U740 ( .A1(n6860), .A2(\mem[163][13] ), .B1(n6828), .B2(
        \mem[184][13] ), .ZN(n405) );
  AOI22D0 U741 ( .A1(n6165), .A2(\mem[174][13] ), .B1(n6748), .B2(
        \mem[169][13] ), .ZN(n404) );
  AOI22D0 U742 ( .A1(n6868), .A2(\mem[171][13] ), .B1(n6760), .B2(
        \mem[173][13] ), .ZN(n402) );
  ND4D0 U743 ( .A1(n405), .A2(n404), .A3(n403), .A4(n402), .ZN(n406) );
  NR4D0 U744 ( .A1(n409), .A2(n408), .A3(n407), .A4(n406), .ZN(n431) );
  AOI22D0 U745 ( .A1(n6903), .A2(\mem[179][13] ), .B1(n6957), .B2(
        \mem[185][13] ), .ZN(n413) );
  AOI22D0 U746 ( .A1(n6928), .A2(\mem[135][13] ), .B1(n6889), .B2(
        \mem[156][13] ), .ZN(n412) );
  AOI22D0 U747 ( .A1(n6923), .A2(\mem[162][13] ), .B1(n6964), .B2(
        \mem[158][13] ), .ZN(n411) );
  AOI22D0 U748 ( .A1(n6914), .A2(\mem[133][13] ), .B1(n6988), .B2(
        \mem[191][13] ), .ZN(n410) );
  ND4D0 U749 ( .A1(n413), .A2(n412), .A3(n411), .A4(n410), .ZN(n429) );
  AOI22D0 U750 ( .A1(n6994), .A2(\mem[190][13] ), .B1(n6804), .B2(
        \mem[147][13] ), .ZN(n417) );
  AOI22D0 U751 ( .A1(n6924), .A2(\mem[160][13] ), .B1(n6906), .B2(
        \mem[140][13] ), .ZN(n416) );
  AOI22D0 U752 ( .A1(n6614), .A2(\mem[150][13] ), .B1(n6174), .B2(
        \mem[182][13] ), .ZN(n415) );
  AOI22D0 U753 ( .A1(n6926), .A2(\mem[129][13] ), .B1(n6847), .B2(
        \mem[153][13] ), .ZN(n414) );
  ND4D0 U754 ( .A1(n417), .A2(n416), .A3(n415), .A4(n414), .ZN(n428) );
  AOI22D0 U755 ( .A1(n6892), .A2(\mem[172][13] ), .B1(n6881), .B2(
        \mem[144][13] ), .ZN(n421) );
  AOI22D0 U756 ( .A1(n6829), .A2(\mem[166][13] ), .B1(n6835), .B2(
        \mem[132][13] ), .ZN(n420) );
  BUFFD0 U757 ( .I(n6888), .Z(n6448) );
  AOI22D0 U758 ( .A1(n6448), .A2(\mem[128][13] ), .B1(n6913), .B2(
        \mem[155][13] ), .ZN(n419) );
  AOI22D0 U759 ( .A1(n6842), .A2(\mem[154][13] ), .B1(n6874), .B2(
        \mem[170][13] ), .ZN(n418) );
  ND4D0 U760 ( .A1(n421), .A2(n420), .A3(n419), .A4(n418), .ZN(n427) );
  AOI22D0 U761 ( .A1(n6959), .A2(\mem[131][13] ), .B1(n6979), .B2(
        \mem[142][13] ), .ZN(n425) );
  AOI22D0 U762 ( .A1(n6728), .A2(\mem[180][13] ), .B1(n6965), .B2(
        \mem[141][13] ), .ZN(n423) );
  AOI22D0 U763 ( .A1(n6659), .A2(\mem[181][13] ), .B1(n6966), .B2(
        \mem[178][13] ), .ZN(n422) );
  NR4D0 U764 ( .A1(n429), .A2(n428), .A3(n427), .A4(n426), .ZN(n430) );
  CKND2D0 U765 ( .A1(n431), .A2(n430), .ZN(n518) );
  AOI22D0 U766 ( .A1(n6883), .A2(\mem[48][13] ), .B1(n6913), .B2(\mem[27][13] ), .ZN(n435) );
  AOI22D0 U767 ( .A1(n6903), .A2(\mem[51][13] ), .B1(n6728), .B2(\mem[52][13] ), .ZN(n434) );
  AOI22D0 U768 ( .A1(n6802), .A2(\mem[24][13] ), .B1(n6698), .B2(\mem[2][13] ), 
        .ZN(n433) );
  AOI22D0 U769 ( .A1(n6933), .A2(\mem[33][13] ), .B1(n6916), .B2(\mem[21][13] ), .ZN(n432) );
  ND4D0 U770 ( .A1(n435), .A2(n434), .A3(n433), .A4(n432), .ZN(n451) );
  AOI22D0 U771 ( .A1(n6873), .A2(\mem[30][13] ), .B1(n6992), .B2(\mem[54][13] ), .ZN(n439) );
  AOI22D0 U772 ( .A1(n6970), .A2(\mem[16][13] ), .B1(n6738), .B2(\mem[37][13] ), .ZN(n438) );
  AOI22D0 U773 ( .A1(n6892), .A2(\mem[44][13] ), .B1(n6733), .B2(\mem[58][13] ), .ZN(n437) );
  AOI22D0 U774 ( .A1(n6907), .A2(\mem[3][13] ), .B1(n6968), .B2(\mem[41][13] ), 
        .ZN(n436) );
  ND4D0 U775 ( .A1(n439), .A2(n438), .A3(n437), .A4(n436), .ZN(n450) );
  AOI22D0 U776 ( .A1(n6868), .A2(\mem[43][13] ), .B1(n6988), .B2(\mem[63][13] ), .ZN(n443) );
  AOI22D0 U777 ( .A1(n6917), .A2(\mem[46][13] ), .B1(n5966), .B2(\mem[31][13] ), .ZN(n442) );
  AOI22D0 U778 ( .A1(n6905), .A2(\mem[59][13] ), .B1(n6842), .B2(\mem[26][13] ), .ZN(n441) );
  AOI22D0 U779 ( .A1(n6747), .A2(\mem[20][13] ), .B1(n6836), .B2(\mem[10][13] ), .ZN(n440) );
  ND4D0 U780 ( .A1(n443), .A2(n442), .A3(n441), .A4(n440), .ZN(n449) );
  AOI22D0 U781 ( .A1(n6993), .A2(\mem[53][13] ), .B1(n6882), .B2(\mem[15][13] ), .ZN(n446) );
  AOI22D0 U782 ( .A1(n6829), .A2(\mem[38][13] ), .B1(n6957), .B2(\mem[57][13] ), .ZN(n445) );
  AOI22D0 U783 ( .A1(n6967), .A2(\mem[39][13] ), .B1(n6809), .B2(\mem[9][13] ), 
        .ZN(n444) );
  ND4D0 U784 ( .A1(n447), .A2(n446), .A3(n445), .A4(n444), .ZN(n448) );
  NR4D0 U785 ( .A1(n451), .A2(n450), .A3(n449), .A4(n448), .ZN(n473) );
  AOI22D0 U786 ( .A1(n6989), .A2(\mem[6][13] ), .B1(n6860), .B2(\mem[35][13] ), 
        .ZN(n455) );
  AOI22D0 U787 ( .A1(n6922), .A2(\mem[29][13] ), .B1(n6906), .B2(\mem[12][13] ), .ZN(n454) );
  AOI22D0 U788 ( .A1(n6870), .A2(\mem[60][13] ), .B1(n6979), .B2(\mem[14][13] ), .ZN(n453) );
  AOI22D0 U789 ( .A1(n6928), .A2(\mem[7][13] ), .B1(n6760), .B2(\mem[45][13] ), 
        .ZN(n452) );
  ND4D0 U790 ( .A1(n455), .A2(n454), .A3(n453), .A4(n452), .ZN(n471) );
  AOI22D0 U791 ( .A1(n6890), .A2(\mem[36][13] ), .B1(n6980), .B2(\mem[61][13] ), .ZN(n459) );
  AOI22D0 U792 ( .A1(n6952), .A2(\mem[22][13] ), .B1(n6814), .B2(\mem[1][13] ), 
        .ZN(n458) );
  AOI22D0 U793 ( .A1(n6880), .A2(\mem[11][13] ), .B1(n6978), .B2(\mem[8][13] ), 
        .ZN(n457) );
  AOI22D0 U794 ( .A1(n6179), .A2(\mem[47][13] ), .B1(n6888), .B2(\mem[0][13] ), 
        .ZN(n456) );
  ND4D0 U795 ( .A1(n459), .A2(n458), .A3(n457), .A4(n456), .ZN(n470) );
  AOI22D0 U796 ( .A1(n6727), .A2(\mem[42][13] ), .B1(n6707), .B2(\mem[23][13] ), .ZN(n463) );
  AOI22D0 U797 ( .A1(n6994), .A2(\mem[62][13] ), .B1(n6658), .B2(\mem[50][13] ), .ZN(n462) );
  AOI22D0 U798 ( .A1(n6923), .A2(\mem[34][13] ), .B1(n6791), .B2(\mem[32][13] ), .ZN(n461) );
  ND4D0 U799 ( .A1(n463), .A2(n462), .A3(n461), .A4(n460), .ZN(n469) );
  AOI22D0 U800 ( .A1(n6956), .A2(\mem[40][13] ), .B1(n6828), .B2(\mem[56][13] ), .ZN(n467) );
  AOI22D0 U801 ( .A1(n6542), .A2(\mem[18][13] ), .B1(n6863), .B2(\mem[55][13] ), .ZN(n466) );
  AOI22D0 U802 ( .A1(n6784), .A2(\mem[28][13] ), .B1(n6904), .B2(\mem[19][13] ), .ZN(n465) );
  AOI22D0 U803 ( .A1(n6835), .A2(\mem[4][13] ), .B1(n6965), .B2(\mem[13][13] ), 
        .ZN(n464) );
  ND4D0 U804 ( .A1(n467), .A2(n466), .A3(n465), .A4(n464), .ZN(n468) );
  NR4D0 U805 ( .A1(n471), .A2(n470), .A3(n469), .A4(n468), .ZN(n472) );
  AOI21D0 U806 ( .A1(n473), .A2(n472), .B(n6856), .ZN(n517) );
  AOI22D0 U807 ( .A1(n6872), .A2(\mem[198][13] ), .B1(n6733), .B2(
        \mem[250][13] ), .ZN(n477) );
  AOI22D0 U808 ( .A1(n6967), .A2(\mem[231][13] ), .B1(n6913), .B2(
        \mem[219][13] ), .ZN(n476) );
  AOI22D0 U809 ( .A1(n6847), .A2(\mem[217][13] ), .B1(n6804), .B2(
        \mem[211][13] ), .ZN(n475) );
  AOI22D0 U810 ( .A1(n6959), .A2(\mem[195][13] ), .B1(n6835), .B2(
        \mem[196][13] ), .ZN(n474) );
  ND4D0 U811 ( .A1(n477), .A2(n476), .A3(n475), .A4(n474), .ZN(n493) );
  AOI22D0 U812 ( .A1(n6814), .A2(\mem[193][13] ), .B1(n6922), .B2(
        \mem[221][13] ), .ZN(n481) );
  AOI22D0 U813 ( .A1(n6915), .A2(\mem[205][13] ), .B1(n6774), .B2(
        \mem[241][13] ), .ZN(n480) );
  AOI22D0 U814 ( .A1(n6883), .A2(\mem[240][13] ), .B1(n6738), .B2(
        \mem[229][13] ), .ZN(n479) );
  AOI22D0 U815 ( .A1(n6890), .A2(\mem[228][13] ), .B1(n6868), .B2(
        \mem[235][13] ), .ZN(n478) );
  ND4D0 U816 ( .A1(n481), .A2(n480), .A3(n479), .A4(n478), .ZN(n492) );
  AOI22D0 U817 ( .A1(n6980), .A2(\mem[253][13] ), .B1(n6952), .B2(
        \mem[214][13] ), .ZN(n485) );
  AOI22D0 U818 ( .A1(n6982), .A2(\mem[194][13] ), .B1(n6978), .B2(
        \mem[200][13] ), .ZN(n484) );
  AOI22D0 U819 ( .A1(n6775), .A2(\mem[236][13] ), .B1(n6988), .B2(
        \mem[255][13] ), .ZN(n482) );
  ND4D0 U820 ( .A1(n485), .A2(n484), .A3(n483), .A4(n482), .ZN(n491) );
  AOI22D0 U821 ( .A1(n6784), .A2(\mem[220][13] ), .B1(n6993), .B2(
        \mem[245][13] ), .ZN(n489) );
  AOI22D0 U822 ( .A1(n6933), .A2(\mem[225][13] ), .B1(n6956), .B2(
        \mem[232][13] ), .ZN(n488) );
  AOI22D0 U823 ( .A1(n6747), .A2(\mem[212][13] ), .B1(n6791), .B2(
        \mem[224][13] ), .ZN(n487) );
  AOI22D0 U824 ( .A1(n6928), .A2(\mem[199][13] ), .B1(n6964), .B2(
        \mem[222][13] ), .ZN(n486) );
  ND4D0 U825 ( .A1(n489), .A2(n488), .A3(n487), .A4(n486), .ZN(n490) );
  NR4D0 U826 ( .A1(n493), .A2(n492), .A3(n491), .A4(n490), .ZN(n515) );
  AOI22D0 U827 ( .A1(n6966), .A2(\mem[242][13] ), .B1(n6836), .B2(
        \mem[202][13] ), .ZN(n497) );
  AOI22D0 U828 ( .A1(n6680), .A2(\mem[223][13] ), .B1(n6992), .B2(
        \mem[246][13] ), .ZN(n496) );
  AOI22D0 U829 ( .A1(n6727), .A2(\mem[234][13] ), .B1(n6936), .B2(
        \mem[209][13] ), .ZN(n495) );
  AOI22D0 U830 ( .A1(n6803), .A2(\mem[247][13] ), .B1(n6901), .B2(
        \mem[201][13] ), .ZN(n494) );
  ND4D0 U831 ( .A1(n497), .A2(n496), .A3(n495), .A4(n494), .ZN(n513) );
  AOI22D0 U832 ( .A1(n6923), .A2(\mem[226][13] ), .B1(n6916), .B2(
        \mem[213][13] ), .ZN(n501) );
  AOI22D0 U833 ( .A1(n6870), .A2(\mem[252][13] ), .B1(n6707), .B2(
        \mem[215][13] ), .ZN(n500) );
  AOI22D0 U834 ( .A1(n6880), .A2(\mem[203][13] ), .B1(n6829), .B2(
        \mem[230][13] ), .ZN(n499) );
  AOI22D0 U835 ( .A1(n6860), .A2(\mem[227][13] ), .B1(n6491), .B2(
        \mem[243][13] ), .ZN(n498) );
  ND4D0 U836 ( .A1(n501), .A2(n500), .A3(n499), .A4(n498), .ZN(n512) );
  AOI22D0 U837 ( .A1(n6530), .A2(\mem[251][13] ), .B1(n6957), .B2(
        \mem[249][13] ), .ZN(n505) );
  AOI22D0 U838 ( .A1(n6759), .A2(\mem[206][13] ), .B1(n6969), .B2(
        \mem[210][13] ), .ZN(n503) );
  AOI22D0 U839 ( .A1(n6917), .A2(\mem[238][13] ), .B1(n6828), .B2(
        \mem[248][13] ), .ZN(n502) );
  AOI22D0 U840 ( .A1(n6953), .A2(\mem[239][13] ), .B1(n6882), .B2(
        \mem[207][13] ), .ZN(n509) );
  AOI22D0 U841 ( .A1(n6934), .A2(\mem[216][13] ), .B1(n6728), .B2(
        \mem[244][13] ), .ZN(n508) );
  AOI22D0 U842 ( .A1(n6754), .A2(\mem[197][13] ), .B1(n6760), .B2(
        \mem[237][13] ), .ZN(n507) );
  AOI22D0 U843 ( .A1(n6881), .A2(\mem[208][13] ), .B1(n6789), .B2(
        \mem[254][13] ), .ZN(n506) );
  ND4D0 U844 ( .A1(n509), .A2(n508), .A3(n507), .A4(n506), .ZN(n510) );
  NR4D0 U845 ( .A1(n513), .A2(n512), .A3(n511), .A4(n510), .ZN(n514) );
  AOI21D0 U846 ( .A1(n515), .A2(n514), .B(n6945), .ZN(n516) );
  AOI211D0 U847 ( .A1(n6951), .A2(n518), .B(n517), .C(n516), .ZN(n540) );
  AOI22D0 U848 ( .A1(n6933), .A2(\mem[97][13] ), .B1(n6993), .B2(
        \mem[117][13] ), .ZN(n522) );
  AOI22D0 U849 ( .A1(n6913), .A2(\mem[91][13] ), .B1(n6956), .B2(
        \mem[104][13] ), .ZN(n521) );
  AOI22D0 U850 ( .A1(n6775), .A2(\mem[108][13] ), .B1(n6967), .B2(
        \mem[103][13] ), .ZN(n520) );
  AOI22D0 U851 ( .A1(n6995), .A2(\mem[87][13] ), .B1(n6738), .B2(
        \mem[101][13] ), .ZN(n519) );
  ND4D0 U852 ( .A1(n522), .A2(n521), .A3(n520), .A4(n519), .ZN(n538) );
  AOI22D0 U853 ( .A1(n6952), .A2(\mem[86][13] ), .B1(n6842), .B2(\mem[90][13] ), .ZN(n526) );
  AOI22D0 U854 ( .A1(n6814), .A2(\mem[65][13] ), .B1(n6906), .B2(\mem[76][13] ), .ZN(n525) );
  AOI22D0 U855 ( .A1(n6733), .A2(\mem[122][13] ), .B1(n6978), .B2(
        \mem[72][13] ), .ZN(n524) );
  ND4D0 U856 ( .A1(n526), .A2(n525), .A3(n524), .A4(n523), .ZN(n537) );
  AOI22D0 U857 ( .A1(n6847), .A2(\mem[89][13] ), .B1(n6958), .B2(\mem[81][13] ), .ZN(n530) );
  AOI22D0 U858 ( .A1(n6870), .A2(\mem[124][13] ), .B1(n6698), .B2(
        \mem[66][13] ), .ZN(n529) );
  AOI22D0 U859 ( .A1(n6861), .A2(\mem[68][13] ), .B1(n6754), .B2(\mem[69][13] ), .ZN(n528) );
  AOI22D0 U860 ( .A1(n6955), .A2(\mem[85][13] ), .B1(n6760), .B2(
        \mem[109][13] ), .ZN(n527) );
  ND4D0 U861 ( .A1(n530), .A2(n529), .A3(n528), .A4(n527), .ZN(n536) );
  AOI22D0 U862 ( .A1(n6928), .A2(\mem[71][13] ), .B1(n6959), .B2(\mem[67][13] ), .ZN(n534) );
  AOI22D0 U863 ( .A1(n6953), .A2(\mem[111][13] ), .B1(n6988), .B2(
        \mem[127][13] ), .ZN(n533) );
  AOI22D0 U864 ( .A1(n6904), .A2(\mem[83][13] ), .B1(n6957), .B2(
        \mem[121][13] ), .ZN(n532) );
  AOI22D0 U865 ( .A1(n6905), .A2(\mem[123][13] ), .B1(n6880), .B2(
        \mem[75][13] ), .ZN(n531) );
  ND4D0 U866 ( .A1(n534), .A2(n533), .A3(n532), .A4(n531), .ZN(n535) );
  NR4D0 U867 ( .A1(n538), .A2(n537), .A3(n536), .A4(n535), .ZN(n539) );
  AOI32D0 U868 ( .A1(n541), .A2(n540), .A3(n539), .B1(n7004), .B2(n540), .ZN(
        dout[13]) );
  AOI22D0 U869 ( .A1(n6995), .A2(\mem[151][15] ), .B1(n6859), .B2(
        \mem[180][15] ), .ZN(n545) );
  AOI22D0 U870 ( .A1(n6966), .A2(\mem[178][15] ), .B1(n6804), .B2(
        \mem[147][15] ), .ZN(n543) );
  AOI22D0 U871 ( .A1(n6958), .A2(\mem[145][15] ), .B1(n6789), .B2(
        \mem[190][15] ), .ZN(n542) );
  ND4D0 U872 ( .A1(n545), .A2(n544), .A3(n543), .A4(n542), .ZN(n561) );
  AOI22D0 U873 ( .A1(n6913), .A2(\mem[155][15] ), .B1(n6680), .B2(
        \mem[159][15] ), .ZN(n549) );
  AOI22D0 U874 ( .A1(n6874), .A2(\mem[170][15] ), .B1(n6976), .B2(
        \mem[162][15] ), .ZN(n548) );
  AOI22D0 U875 ( .A1(n6922), .A2(\mem[157][15] ), .B1(n6659), .B2(
        \mem[181][15] ), .ZN(n547) );
  AOI22D0 U876 ( .A1(n6903), .A2(\mem[179][15] ), .B1(n6927), .B2(
        \mem[153][15] ), .ZN(n546) );
  ND4D0 U877 ( .A1(n549), .A2(n548), .A3(n547), .A4(n546), .ZN(n560) );
  AOI22D0 U878 ( .A1(n6837), .A2(\mem[143][15] ), .B1(n6964), .B2(
        \mem[158][15] ), .ZN(n553) );
  AOI22D0 U879 ( .A1(n6563), .A2(\mem[136][15] ), .B1(n6902), .B2(
        \mem[165][15] ), .ZN(n552) );
  AOI22D0 U880 ( .A1(n6869), .A2(\mem[177][15] ), .B1(n6174), .B2(
        \mem[182][15] ), .ZN(n551) );
  AOI22D0 U881 ( .A1(n6828), .A2(\mem[184][15] ), .B1(n6990), .B2(
        \mem[140][15] ), .ZN(n550) );
  ND4D0 U882 ( .A1(n553), .A2(n552), .A3(n551), .A4(n550), .ZN(n559) );
  AOI22D0 U883 ( .A1(n6982), .A2(\mem[130][15] ), .B1(n6748), .B2(
        \mem[169][15] ), .ZN(n557) );
  AOI22D0 U884 ( .A1(n6954), .A2(\mem[138][15] ), .B1(n6935), .B2(
        \mem[191][15] ), .ZN(n556) );
  AOI22D0 U885 ( .A1(n6915), .A2(\mem[141][15] ), .B1(n6925), .B2(
        \mem[173][15] ), .ZN(n555) );
  ND4D0 U886 ( .A1(n557), .A2(n556), .A3(n555), .A4(n554), .ZN(n558) );
  NR4D0 U887 ( .A1(n561), .A2(n560), .A3(n559), .A4(n558), .ZN(n4809) );
  INVD0 U888 ( .I(n7004), .ZN(n6164) );
  AOI22D0 U889 ( .A1(n6784), .A2(\mem[92][15] ), .B1(n6869), .B2(
        \mem[113][15] ), .ZN(n565) );
  AOI22D0 U890 ( .A1(n6923), .A2(\mem[98][15] ), .B1(n6760), .B2(
        \mem[109][15] ), .ZN(n564) );
  AOI22D0 U891 ( .A1(n6775), .A2(\mem[108][15] ), .B1(n6871), .B2(
        \mem[121][15] ), .ZN(n563) );
  AOI22D0 U892 ( .A1(n6967), .A2(\mem[103][15] ), .B1(n6956), .B2(
        \mem[104][15] ), .ZN(n562) );
  ND4D0 U893 ( .A1(n565), .A2(n564), .A3(n563), .A4(n562), .ZN(n4677) );
  AOI22D0 U894 ( .A1(n6179), .A2(\mem[111][15] ), .B1(n6802), .B2(
        \mem[88][15] ), .ZN(n569) );
  AOI22D0 U895 ( .A1(n6981), .A2(\mem[124][15] ), .B1(n6964), .B2(
        \mem[94][15] ), .ZN(n568) );
  AOI22D0 U896 ( .A1(n6819), .A2(\mem[125][15] ), .B1(n6906), .B2(
        \mem[76][15] ), .ZN(n566) );
  ND4D0 U897 ( .A1(n569), .A2(n568), .A3(n567), .A4(n566), .ZN(n4676) );
  AOI22D0 U898 ( .A1(n6971), .A2(\mem[102][15] ), .B1(n6863), .B2(
        \mem[119][15] ), .ZN(n4669) );
  AOI22D0 U899 ( .A1(n6969), .A2(\mem[82][15] ), .B1(n6988), .B2(
        \mem[127][15] ), .ZN(n572) );
  AOI22D0 U900 ( .A1(n6883), .A2(\mem[112][15] ), .B1(n6992), .B2(
        \mem[118][15] ), .ZN(n571) );
  AOI22D0 U901 ( .A1(n6847), .A2(\mem[89][15] ), .B1(n6966), .B2(
        \mem[114][15] ), .ZN(n570) );
  ND4D0 U902 ( .A1(n4669), .A2(n572), .A3(n571), .A4(n570), .ZN(n4675) );
  AOI22D0 U903 ( .A1(n6830), .A2(\mem[71][15] ), .B1(n6952), .B2(\mem[86][15] ), .ZN(n4673) );
  AOI22D0 U904 ( .A1(n6814), .A2(\mem[65][15] ), .B1(n6491), .B2(
        \mem[115][15] ), .ZN(n4672) );
  AOI22D0 U905 ( .A1(n6888), .A2(\mem[64][15] ), .B1(n6936), .B2(\mem[81][15] ), .ZN(n4671) );
  AOI22D0 U906 ( .A1(n6861), .A2(\mem[68][15] ), .B1(n6842), .B2(\mem[90][15] ), .ZN(n4670) );
  ND4D0 U907 ( .A1(n4673), .A2(n4672), .A3(n4671), .A4(n4670), .ZN(n4674) );
  NR4D0 U908 ( .A1(n4677), .A2(n4676), .A3(n4675), .A4(n4674), .ZN(n4699) );
  AOI22D0 U909 ( .A1(n6978), .A2(\mem[72][15] ), .B1(n6912), .B2(
        \mem[120][15] ), .ZN(n4681) );
  AOI22D0 U910 ( .A1(n6955), .A2(\mem[85][15] ), .B1(n6837), .B2(\mem[79][15] ), .ZN(n4680) );
  AOI22D0 U911 ( .A1(n6933), .A2(\mem[97][15] ), .B1(n6879), .B2(
        \mem[122][15] ), .ZN(n4679) );
  AOI22D0 U912 ( .A1(n6970), .A2(\mem[80][15] ), .B1(n6904), .B2(\mem[83][15] ), .ZN(n4678) );
  ND4D0 U913 ( .A1(n4681), .A2(n4680), .A3(n4679), .A4(n4678), .ZN(n4697) );
  AOI22D0 U914 ( .A1(n6880), .A2(\mem[75][15] ), .B1(n6754), .B2(\mem[69][15] ), .ZN(n4685) );
  AOI22D0 U915 ( .A1(n6872), .A2(\mem[70][15] ), .B1(n6698), .B2(\mem[66][15] ), .ZN(n4683) );
  AOI22D0 U916 ( .A1(n6913), .A2(\mem[91][15] ), .B1(n6748), .B2(
        \mem[105][15] ), .ZN(n4682) );
  ND4D0 U917 ( .A1(n4685), .A2(n4684), .A3(n4683), .A4(n4682), .ZN(n4696) );
  AOI22D0 U918 ( .A1(n6525), .A2(\mem[99][15] ), .B1(n6954), .B2(\mem[74][15] ), .ZN(n4689) );
  AOI22D0 U919 ( .A1(n6901), .A2(\mem[73][15] ), .B1(n6738), .B2(
        \mem[101][15] ), .ZN(n4688) );
  AOI22D0 U920 ( .A1(n6165), .A2(\mem[110][15] ), .B1(n6915), .B2(
        \mem[77][15] ), .ZN(n4687) );
  AOI22D0 U921 ( .A1(n6759), .A2(\mem[78][15] ), .B1(n6868), .B2(
        \mem[107][15] ), .ZN(n4686) );
  ND4D0 U922 ( .A1(n4689), .A2(n4688), .A3(n4687), .A4(n4686), .ZN(n4695) );
  AOI22D0 U923 ( .A1(n6907), .A2(\mem[67][15] ), .B1(n6995), .B2(\mem[87][15] ), .ZN(n4693) );
  AOI22D0 U924 ( .A1(n6922), .A2(\mem[93][15] ), .B1(n6993), .B2(
        \mem[117][15] ), .ZN(n4692) );
  AOI22D0 U925 ( .A1(n6680), .A2(\mem[95][15] ), .B1(n6791), .B2(\mem[96][15] ), .ZN(n4691) );
  AOI22D0 U926 ( .A1(n6773), .A2(\mem[100][15] ), .B1(n6789), .B2(
        \mem[126][15] ), .ZN(n4690) );
  ND4D0 U927 ( .A1(n4693), .A2(n4692), .A3(n4691), .A4(n4690), .ZN(n4694) );
  NR4D0 U928 ( .A1(n4697), .A2(n4696), .A3(n4695), .A4(n4694), .ZN(n4698) );
  CKND2D0 U929 ( .A1(n4699), .A2(n4698), .ZN(n4786) );
  AOI22D0 U930 ( .A1(n6847), .A2(\mem[217][15] ), .B1(n6988), .B2(
        \mem[255][15] ), .ZN(n4703) );
  AOI22D0 U931 ( .A1(n6868), .A2(\mem[235][15] ), .B1(n6904), .B2(
        \mem[211][15] ), .ZN(n4702) );
  AOI22D0 U932 ( .A1(n6953), .A2(\mem[239][15] ), .B1(n6923), .B2(
        \mem[226][15] ), .ZN(n4701) );
  AOI22D0 U933 ( .A1(n6530), .A2(\mem[251][15] ), .B1(n6922), .B2(
        \mem[221][15] ), .ZN(n4700) );
  AOI22D0 U934 ( .A1(n6891), .A2(\mem[218][15] ), .B1(n6760), .B2(
        \mem[237][15] ), .ZN(n4706) );
  AOI22D0 U935 ( .A1(n6914), .A2(\mem[197][15] ), .B1(n6874), .B2(
        \mem[234][15] ), .ZN(n4705) );
  AOI22D0 U936 ( .A1(n6759), .A2(\mem[206][15] ), .B1(n6992), .B2(
        \mem[246][15] ), .ZN(n4704) );
  ND4D0 U937 ( .A1(n4707), .A2(n4706), .A3(n4705), .A4(n4704), .ZN(n4718) );
  AOI22D0 U938 ( .A1(n6967), .A2(\mem[231][15] ), .B1(n6916), .B2(
        \mem[213][15] ), .ZN(n4711) );
  AOI22D0 U939 ( .A1(n6809), .A2(\mem[201][15] ), .B1(n6936), .B2(
        \mem[209][15] ), .ZN(n4710) );
  AOI22D0 U940 ( .A1(n6525), .A2(\mem[227][15] ), .B1(n6956), .B2(
        \mem[232][15] ), .ZN(n4709) );
  AOI22D0 U941 ( .A1(n6934), .A2(\mem[216][15] ), .B1(n6913), .B2(
        \mem[219][15] ), .ZN(n4708) );
  ND4D0 U942 ( .A1(n4711), .A2(n4710), .A3(n4709), .A4(n4708), .ZN(n4717) );
  AOI22D0 U943 ( .A1(n6971), .A2(\mem[230][15] ), .B1(n6836), .B2(
        \mem[202][15] ), .ZN(n4715) );
  AOI22D0 U944 ( .A1(n5966), .A2(\mem[223][15] ), .B1(n6964), .B2(
        \mem[222][15] ), .ZN(n4714) );
  AOI22D0 U945 ( .A1(n6448), .A2(\mem[192][15] ), .B1(n6491), .B2(
        \mem[243][15] ), .ZN(n4713) );
  AOI22D0 U946 ( .A1(n6933), .A2(\mem[225][15] ), .B1(n6879), .B2(
        \mem[250][15] ), .ZN(n4712) );
  ND4D0 U947 ( .A1(n4715), .A2(n4714), .A3(n4713), .A4(n4712), .ZN(n4716) );
  NR4D0 U948 ( .A1(n4719), .A2(n4718), .A3(n4717), .A4(n4716), .ZN(n4741) );
  AOI22D0 U949 ( .A1(n6883), .A2(\mem[240][15] ), .B1(n6748), .B2(
        \mem[233][15] ), .ZN(n4723) );
  AOI22D0 U950 ( .A1(n6889), .A2(\mem[220][15] ), .B1(n6728), .B2(
        \mem[244][15] ), .ZN(n4722) );
  AOI22D0 U951 ( .A1(n6981), .A2(\mem[252][15] ), .B1(n6993), .B2(
        \mem[245][15] ), .ZN(n4721) );
  ND4D0 U952 ( .A1(n4723), .A2(n4722), .A3(n4721), .A4(n4720), .ZN(n4739) );
  AOI22D0 U953 ( .A1(n6863), .A2(\mem[247][15] ), .B1(n6563), .B2(
        \mem[200][15] ), .ZN(n4727) );
  AOI22D0 U954 ( .A1(n6892), .A2(\mem[236][15] ), .B1(n6989), .B2(
        \mem[198][15] ), .ZN(n4726) );
  AOI22D0 U955 ( .A1(n6970), .A2(\mem[208][15] ), .B1(n6966), .B2(
        \mem[242][15] ), .ZN(n4725) );
  AOI22D0 U956 ( .A1(n6952), .A2(\mem[214][15] ), .B1(n6707), .B2(
        \mem[215][15] ), .ZN(n4724) );
  ND4D0 U957 ( .A1(n4727), .A2(n4726), .A3(n4725), .A4(n4724), .ZN(n4738) );
  AOI22D0 U958 ( .A1(n6917), .A2(\mem[238][15] ), .B1(n6738), .B2(
        \mem[229][15] ), .ZN(n4731) );
  AOI22D0 U959 ( .A1(n6890), .A2(\mem[228][15] ), .B1(n6791), .B2(
        \mem[224][15] ), .ZN(n4730) );
  AOI22D0 U960 ( .A1(n6819), .A2(\mem[253][15] ), .B1(n6959), .B2(
        \mem[195][15] ), .ZN(n4729) );
  AOI22D0 U961 ( .A1(n6928), .A2(\mem[199][15] ), .B1(n6835), .B2(
        \mem[196][15] ), .ZN(n4728) );
  ND4D0 U962 ( .A1(n4731), .A2(n4730), .A3(n4729), .A4(n4728), .ZN(n4737) );
  AOI22D0 U963 ( .A1(n6926), .A2(\mem[193][15] ), .B1(n6698), .B2(
        \mem[194][15] ), .ZN(n4735) );
  AOI22D0 U964 ( .A1(n6965), .A2(\mem[205][15] ), .B1(n6882), .B2(
        \mem[207][15] ), .ZN(n4734) );
  AOI22D0 U965 ( .A1(n6542), .A2(\mem[210][15] ), .B1(n6774), .B2(
        \mem[241][15] ), .ZN(n4733) );
  AOI22D0 U966 ( .A1(n6325), .A2(\mem[203][15] ), .B1(n6828), .B2(
        \mem[248][15] ), .ZN(n4732) );
  ND4D0 U967 ( .A1(n4735), .A2(n4734), .A3(n4733), .A4(n4732), .ZN(n4736) );
  NR4D0 U968 ( .A1(n4739), .A2(n4738), .A3(n4737), .A4(n4736), .ZN(n4740) );
  AOI21D0 U969 ( .A1(n4741), .A2(n4740), .B(n6945), .ZN(n4785) );
  AOI22D0 U970 ( .A1(n6993), .A2(\mem[53][15] ), .B1(n6978), .B2(\mem[8][15] ), 
        .ZN(n4745) );
  AOI22D0 U971 ( .A1(n6913), .A2(\mem[27][15] ), .B1(n6707), .B2(\mem[23][15] ), .ZN(n4744) );
  AOI22D0 U972 ( .A1(n6879), .A2(\mem[58][15] ), .B1(n6847), .B2(\mem[25][15] ), .ZN(n4742) );
  ND4D0 U973 ( .A1(n4745), .A2(n4744), .A3(n4743), .A4(n4742), .ZN(n4761) );
  AOI22D0 U974 ( .A1(n6863), .A2(\mem[55][15] ), .B1(n6874), .B2(\mem[42][15] ), .ZN(n4749) );
  AOI22D0 U975 ( .A1(n6980), .A2(\mem[61][15] ), .B1(n6871), .B2(\mem[57][15] ), .ZN(n4748) );
  AOI22D0 U976 ( .A1(n6889), .A2(\mem[28][15] ), .B1(n6728), .B2(\mem[52][15] ), .ZN(n4747) );
  AOI22D0 U977 ( .A1(n6542), .A2(\mem[18][15] ), .B1(n6901), .B2(\mem[9][15] ), 
        .ZN(n4746) );
  ND4D0 U978 ( .A1(n4749), .A2(n4748), .A3(n4747), .A4(n4746), .ZN(n4760) );
  AOI22D0 U979 ( .A1(n6926), .A2(\mem[1][15] ), .B1(n6774), .B2(\mem[49][15] ), 
        .ZN(n4753) );
  AOI22D0 U980 ( .A1(n6953), .A2(\mem[47][15] ), .B1(n6966), .B2(\mem[50][15] ), .ZN(n4752) );
  AOI22D0 U981 ( .A1(n6925), .A2(\mem[45][15] ), .B1(n6738), .B2(\mem[37][15] ), .ZN(n4751) );
  AOI22D0 U982 ( .A1(n6890), .A2(\mem[36][15] ), .B1(n6956), .B2(\mem[40][15] ), .ZN(n4750) );
  ND4D0 U983 ( .A1(n4753), .A2(n4752), .A3(n4751), .A4(n4750), .ZN(n4759) );
  AOI22D0 U984 ( .A1(n6933), .A2(\mem[33][15] ), .B1(n6789), .B2(\mem[62][15] ), .ZN(n4757) );
  AOI22D0 U985 ( .A1(n6959), .A2(\mem[3][15] ), .B1(n6983), .B2(\mem[48][15] ), 
        .ZN(n4756) );
  AOI22D0 U986 ( .A1(n6989), .A2(\mem[6][15] ), .B1(n6860), .B2(\mem[35][15] ), 
        .ZN(n4755) );
  AOI22D0 U987 ( .A1(n6904), .A2(\mem[19][15] ), .B1(n6988), .B2(\mem[63][15] ), .ZN(n4754) );
  ND4D0 U988 ( .A1(n4757), .A2(n4756), .A3(n4755), .A4(n4754), .ZN(n4758) );
  NR4D0 U989 ( .A1(n4761), .A2(n4760), .A3(n4759), .A4(n4758), .ZN(n4783) );
  AOI22D0 U990 ( .A1(n6934), .A2(\mem[24][15] ), .B1(n6828), .B2(\mem[56][15] ), .ZN(n4765) );
  AOI22D0 U991 ( .A1(n6914), .A2(\mem[5][15] ), .B1(n6680), .B2(\mem[31][15] ), 
        .ZN(n4763) );
  AOI22D0 U992 ( .A1(n6979), .A2(\mem[14][15] ), .B1(n6916), .B2(\mem[21][15] ), .ZN(n4762) );
  ND4D0 U993 ( .A1(n4765), .A2(n4764), .A3(n4763), .A4(n4762), .ZN(n4781) );
  AOI22D0 U994 ( .A1(n6970), .A2(\mem[16][15] ), .B1(n6936), .B2(\mem[17][15] ), .ZN(n4769) );
  AOI22D0 U995 ( .A1(n6982), .A2(\mem[2][15] ), .B1(n6882), .B2(\mem[15][15] ), 
        .ZN(n4768) );
  AOI22D0 U996 ( .A1(n6991), .A2(\mem[20][15] ), .B1(n6964), .B2(\mem[30][15] ), .ZN(n4767) );
  AOI22D0 U997 ( .A1(n6917), .A2(\mem[46][15] ), .B1(n6491), .B2(\mem[51][15] ), .ZN(n4766) );
  ND4D0 U998 ( .A1(n4769), .A2(n4768), .A3(n4767), .A4(n4766), .ZN(n4780) );
  AOI22D0 U999 ( .A1(n6928), .A2(\mem[7][15] ), .B1(n6906), .B2(\mem[12][15] ), 
        .ZN(n4773) );
  AOI22D0 U1000 ( .A1(n6880), .A2(\mem[11][15] ), .B1(n6891), .B2(
        \mem[26][15] ), .ZN(n4772) );
  AOI22D0 U1001 ( .A1(n6835), .A2(\mem[4][15] ), .B1(n6639), .B2(\mem[39][15] ), .ZN(n4771) );
  AOI22D0 U1002 ( .A1(n6922), .A2(\mem[29][15] ), .B1(n6174), .B2(
        \mem[54][15] ), .ZN(n4770) );
  ND4D0 U1003 ( .A1(n4773), .A2(n4772), .A3(n4771), .A4(n4770), .ZN(n4779) );
  AOI22D0 U1004 ( .A1(n6829), .A2(\mem[38][15] ), .B1(n6791), .B2(
        \mem[32][15] ), .ZN(n4777) );
  AOI22D0 U1005 ( .A1(n6868), .A2(\mem[43][15] ), .B1(n6888), .B2(\mem[0][15] ), .ZN(n4776) );
  AOI22D0 U1006 ( .A1(n6954), .A2(\mem[10][15] ), .B1(n6965), .B2(
        \mem[13][15] ), .ZN(n4775) );
  AOI22D0 U1007 ( .A1(n6952), .A2(\mem[22][15] ), .B1(n6748), .B2(
        \mem[41][15] ), .ZN(n4774) );
  NR4D0 U1008 ( .A1(n4781), .A2(n4780), .A3(n4779), .A4(n4778), .ZN(n4782) );
  AOI21D0 U1009 ( .A1(n4783), .A2(n4782), .B(n6856), .ZN(n4784) );
  AOI211D0 U1010 ( .A1(n6164), .A2(n4786), .B(n4785), .C(n4784), .ZN(n4808) );
  AOI22D0 U1011 ( .A1(n6892), .A2(\mem[172][15] ), .B1(n6952), .B2(
        \mem[150][15] ), .ZN(n4790) );
  AOI22D0 U1012 ( .A1(n6759), .A2(\mem[142][15] ), .B1(n6868), .B2(
        \mem[171][15] ), .ZN(n4789) );
  AOI22D0 U1013 ( .A1(n6989), .A2(\mem[134][15] ), .B1(n6926), .B2(
        \mem[129][15] ), .ZN(n4788) );
  AOI22D0 U1014 ( .A1(n6905), .A2(\mem[187][15] ), .B1(n6880), .B2(
        \mem[139][15] ), .ZN(n4787) );
  ND4D0 U1015 ( .A1(n4790), .A2(n4789), .A3(n4788), .A4(n4787), .ZN(n4806) );
  AOI22D0 U1016 ( .A1(n6165), .A2(\mem[174][15] ), .B1(n6802), .B2(
        \mem[152][15] ), .ZN(n4794) );
  AOI22D0 U1017 ( .A1(n6179), .A2(\mem[175][15] ), .B1(n6890), .B2(
        \mem[164][15] ), .ZN(n4793) );
  AOI22D0 U1018 ( .A1(n6980), .A2(\mem[189][15] ), .B1(n6959), .B2(
        \mem[131][15] ), .ZN(n4792) );
  AOI22D0 U1019 ( .A1(n6928), .A2(\mem[135][15] ), .B1(n6981), .B2(
        \mem[188][15] ), .ZN(n4791) );
  ND4D0 U1020 ( .A1(n4794), .A2(n4793), .A3(n4792), .A4(n4791), .ZN(n4805) );
  AOI22D0 U1021 ( .A1(n6448), .A2(\mem[128][15] ), .B1(n6863), .B2(
        \mem[183][15] ), .ZN(n4798) );
  AOI22D0 U1022 ( .A1(n6754), .A2(\mem[133][15] ), .B1(n6901), .B2(
        \mem[137][15] ), .ZN(n4796) );
  AOI22D0 U1023 ( .A1(n6733), .A2(\mem[186][15] ), .B1(n6842), .B2(
        \mem[154][15] ), .ZN(n4795) );
  ND4D0 U1024 ( .A1(n4798), .A2(n4797), .A3(n4796), .A4(n4795), .ZN(n4804) );
  AOI22D0 U1025 ( .A1(n6784), .A2(\mem[156][15] ), .B1(n6829), .B2(
        \mem[166][15] ), .ZN(n4802) );
  AOI22D0 U1026 ( .A1(n6747), .A2(\mem[148][15] ), .B1(n6860), .B2(
        \mem[163][15] ), .ZN(n4801) );
  AOI22D0 U1027 ( .A1(n6835), .A2(\mem[132][15] ), .B1(n6639), .B2(
        \mem[167][15] ), .ZN(n4800) );
  AOI22D0 U1028 ( .A1(n6883), .A2(\mem[176][15] ), .B1(n6933), .B2(
        \mem[161][15] ), .ZN(n4799) );
  NR4D0 U1029 ( .A1(n4806), .A2(n4805), .A3(n4804), .A4(n4803), .ZN(n4807) );
  AOI32D0 U1030 ( .A1(n4809), .A2(n4808), .A3(n4807), .B1(n6188), .B2(n4808), 
        .ZN(dout[15]) );
  AOI22D0 U1031 ( .A1(n6727), .A2(\mem[106][14] ), .B1(n6760), .B2(
        \mem[109][14] ), .ZN(n4813) );
  AOI22D0 U1032 ( .A1(n6967), .A2(\mem[103][14] ), .B1(n6836), .B2(
        \mem[74][14] ), .ZN(n4812) );
  AOI22D0 U1033 ( .A1(n6917), .A2(\mem[110][14] ), .B1(n6791), .B2(
        \mem[96][14] ), .ZN(n4811) );
  AOI22D0 U1034 ( .A1(n6904), .A2(\mem[83][14] ), .B1(n6978), .B2(
        \mem[72][14] ), .ZN(n4810) );
  ND4D0 U1035 ( .A1(n4813), .A2(n4812), .A3(n4811), .A4(n4810), .ZN(n4829) );
  AOI22D0 U1036 ( .A1(n6935), .A2(\mem[127][14] ), .B1(n6871), .B2(
        \mem[121][14] ), .ZN(n4817) );
  AOI22D0 U1037 ( .A1(n6870), .A2(\mem[124][14] ), .B1(n6882), .B2(
        \mem[79][14] ), .ZN(n4816) );
  AOI22D0 U1038 ( .A1(n6747), .A2(\mem[84][14] ), .B1(n6992), .B2(
        \mem[118][14] ), .ZN(n4815) );
  AOI22D0 U1039 ( .A1(n6759), .A2(\mem[78][14] ), .B1(n6860), .B2(
        \mem[99][14] ), .ZN(n4814) );
  ND4D0 U1040 ( .A1(n4817), .A2(n4816), .A3(n4815), .A4(n4814), .ZN(n4828) );
  AOI22D0 U1041 ( .A1(n6980), .A2(\mem[125][14] ), .B1(n6901), .B2(
        \mem[73][14] ), .ZN(n4821) );
  AOI22D0 U1042 ( .A1(n6888), .A2(\mem[64][14] ), .B1(n6728), .B2(
        \mem[116][14] ), .ZN(n4819) );
  AOI22D0 U1043 ( .A1(n6754), .A2(\mem[69][14] ), .B1(n6916), .B2(
        \mem[85][14] ), .ZN(n4818) );
  ND4D0 U1044 ( .A1(n4821), .A2(n4820), .A3(n4819), .A4(n4818), .ZN(n4827) );
  AOI22D0 U1045 ( .A1(n6863), .A2(\mem[119][14] ), .B1(n6964), .B2(
        \mem[94][14] ), .ZN(n4825) );
  AOI22D0 U1046 ( .A1(n6883), .A2(\mem[112][14] ), .B1(n6956), .B2(
        \mem[104][14] ), .ZN(n4824) );
  AOI22D0 U1047 ( .A1(n6880), .A2(\mem[75][14] ), .B1(n6989), .B2(
        \mem[70][14] ), .ZN(n4823) );
  AOI22D0 U1048 ( .A1(n6952), .A2(\mem[86][14] ), .B1(n6922), .B2(
        \mem[93][14] ), .ZN(n4822) );
  ND4D0 U1049 ( .A1(n4825), .A2(n4824), .A3(n4823), .A4(n4822), .ZN(n4826) );
  NR4D0 U1050 ( .A1(n4829), .A2(n4828), .A3(n4827), .A4(n4826), .ZN(n4981) );
  AOI22D0 U1051 ( .A1(n6728), .A2(\mem[180][14] ), .B1(n6738), .B2(
        \mem[165][14] ), .ZN(n4833) );
  AOI22D0 U1052 ( .A1(n6847), .A2(\mem[153][14] ), .B1(n6828), .B2(
        \mem[184][14] ), .ZN(n4832) );
  AOI22D0 U1053 ( .A1(n6967), .A2(\mem[167][14] ), .B1(n6901), .B2(
        \mem[137][14] ), .ZN(n4831) );
  AOI22D0 U1054 ( .A1(n6784), .A2(\mem[156][14] ), .B1(n6906), .B2(
        \mem[140][14] ), .ZN(n4830) );
  ND4D0 U1055 ( .A1(n4833), .A2(n4832), .A3(n4831), .A4(n4830), .ZN(n4849) );
  AOI22D0 U1056 ( .A1(n6733), .A2(\mem[186][14] ), .B1(n6789), .B2(
        \mem[190][14] ), .ZN(n4837) );
  AOI22D0 U1057 ( .A1(n6926), .A2(\mem[129][14] ), .B1(n6842), .B2(
        \mem[154][14] ), .ZN(n4836) );
  AOI22D0 U1058 ( .A1(n6964), .A2(\mem[158][14] ), .B1(n6774), .B2(
        \mem[177][14] ), .ZN(n4835) );
  AOI22D0 U1059 ( .A1(n6542), .A2(\mem[146][14] ), .B1(n6874), .B2(
        \mem[170][14] ), .ZN(n4834) );
  ND4D0 U1060 ( .A1(n4837), .A2(n4836), .A3(n4835), .A4(n4834), .ZN(n4848) );
  AOI22D0 U1061 ( .A1(n6959), .A2(\mem[131][14] ), .B1(n6658), .B2(
        \mem[178][14] ), .ZN(n4841) );
  AOI22D0 U1062 ( .A1(n6981), .A2(\mem[188][14] ), .B1(n6882), .B2(
        \mem[143][14] ), .ZN(n4840) );
  AOI22D0 U1063 ( .A1(n6880), .A2(\mem[139][14] ), .B1(n6978), .B2(
        \mem[136][14] ), .ZN(n4839) );
  AOI22D0 U1064 ( .A1(n6892), .A2(\mem[172][14] ), .B1(n6993), .B2(
        \mem[181][14] ), .ZN(n4838) );
  AOI22D0 U1065 ( .A1(n6989), .A2(\mem[134][14] ), .B1(n6913), .B2(
        \mem[155][14] ), .ZN(n4844) );
  AOI22D0 U1066 ( .A1(n6829), .A2(\mem[166][14] ), .B1(n6804), .B2(
        \mem[147][14] ), .ZN(n4843) );
  AOI22D0 U1067 ( .A1(n6988), .A2(\mem[191][14] ), .B1(n6698), .B2(
        \mem[130][14] ), .ZN(n4842) );
  ND4D0 U1068 ( .A1(n4845), .A2(n4844), .A3(n4843), .A4(n4842), .ZN(n4846) );
  NR4D0 U1069 ( .A1(n4849), .A2(n4848), .A3(n4847), .A4(n4846), .ZN(n4871) );
  AOI22D0 U1070 ( .A1(n6917), .A2(\mem[174][14] ), .B1(n6802), .B2(
        \mem[152][14] ), .ZN(n4853) );
  AOI22D0 U1071 ( .A1(n6923), .A2(\mem[162][14] ), .B1(n6956), .B2(
        \mem[168][14] ), .ZN(n4852) );
  AOI22D0 U1072 ( .A1(n6980), .A2(\mem[189][14] ), .B1(n5966), .B2(
        \mem[159][14] ), .ZN(n4851) );
  AOI22D0 U1073 ( .A1(n6914), .A2(\mem[133][14] ), .B1(n6992), .B2(
        \mem[182][14] ), .ZN(n4850) );
  ND4D0 U1074 ( .A1(n4853), .A2(n4852), .A3(n4851), .A4(n4850), .ZN(n4869) );
  AOI22D0 U1075 ( .A1(n6883), .A2(\mem[176][14] ), .B1(n6965), .B2(
        \mem[141][14] ), .ZN(n4857) );
  AOI22D0 U1076 ( .A1(n6868), .A2(\mem[171][14] ), .B1(n6860), .B2(
        \mem[163][14] ), .ZN(n4856) );
  AOI22D0 U1077 ( .A1(n6759), .A2(\mem[142][14] ), .B1(n6936), .B2(
        \mem[145][14] ), .ZN(n4855) );
  AOI22D0 U1078 ( .A1(n6861), .A2(\mem[132][14] ), .B1(n6707), .B2(
        \mem[151][14] ), .ZN(n4854) );
  ND4D0 U1079 ( .A1(n4857), .A2(n4856), .A3(n4855), .A4(n4854), .ZN(n4868) );
  AOI22D0 U1080 ( .A1(n6953), .A2(\mem[175][14] ), .B1(n6836), .B2(
        \mem[138][14] ), .ZN(n4861) );
  AOI22D0 U1081 ( .A1(n6903), .A2(\mem[179][14] ), .B1(n6760), .B2(
        \mem[173][14] ), .ZN(n4860) );
  AOI22D0 U1082 ( .A1(n6614), .A2(\mem[150][14] ), .B1(n6863), .B2(
        \mem[183][14] ), .ZN(n4859) );
  ND4D0 U1083 ( .A1(n4861), .A2(n4860), .A3(n4859), .A4(n4858), .ZN(n4867) );
  AOI22D0 U1084 ( .A1(n6890), .A2(\mem[164][14] ), .B1(n6933), .B2(
        \mem[161][14] ), .ZN(n4865) );
  AOI22D0 U1085 ( .A1(n6881), .A2(\mem[144][14] ), .B1(n6916), .B2(
        \mem[149][14] ), .ZN(n4864) );
  AOI22D0 U1086 ( .A1(n6928), .A2(\mem[135][14] ), .B1(n6922), .B2(
        \mem[157][14] ), .ZN(n4863) );
  AOI22D0 U1087 ( .A1(n6448), .A2(\mem[128][14] ), .B1(n6791), .B2(
        \mem[160][14] ), .ZN(n4862) );
  ND4D0 U1088 ( .A1(n4865), .A2(n4864), .A3(n4863), .A4(n4862), .ZN(n4866) );
  NR4D0 U1089 ( .A1(n4869), .A2(n4868), .A3(n4867), .A4(n4866), .ZN(n4870) );
  CKND2D0 U1090 ( .A1(n4871), .A2(n4870), .ZN(n4958) );
  AOI22D0 U1091 ( .A1(n6749), .A2(\mem[235][14] ), .B1(n6491), .B2(
        \mem[243][14] ), .ZN(n4875) );
  AOI22D0 U1092 ( .A1(n6889), .A2(\mem[220][14] ), .B1(n6993), .B2(
        \mem[245][14] ), .ZN(n4874) );
  AOI22D0 U1093 ( .A1(n6994), .A2(\mem[254][14] ), .B1(n6738), .B2(
        \mem[229][14] ), .ZN(n4873) );
  AOI22D0 U1094 ( .A1(n6835), .A2(\mem[196][14] ), .B1(n6964), .B2(
        \mem[222][14] ), .ZN(n4872) );
  ND4D0 U1095 ( .A1(n4875), .A2(n4874), .A3(n4873), .A4(n4872), .ZN(n4891) );
  AOI22D0 U1096 ( .A1(n6923), .A2(\mem[226][14] ), .B1(n6988), .B2(
        \mem[255][14] ), .ZN(n4879) );
  AOI22D0 U1097 ( .A1(n6953), .A2(\mem[239][14] ), .B1(n6936), .B2(
        \mem[209][14] ), .ZN(n4878) );
  AOI22D0 U1098 ( .A1(n6952), .A2(\mem[214][14] ), .B1(n6698), .B2(
        \mem[194][14] ), .ZN(n4877) );
  AOI22D0 U1099 ( .A1(n6880), .A2(\mem[203][14] ), .B1(n6926), .B2(
        \mem[193][14] ), .ZN(n4876) );
  ND4D0 U1100 ( .A1(n4879), .A2(n4878), .A3(n4877), .A4(n4876), .ZN(n4890) );
  AOI22D0 U1101 ( .A1(n6959), .A2(\mem[195][14] ), .B1(n6881), .B2(
        \mem[208][14] ), .ZN(n4883) );
  AOI22D0 U1102 ( .A1(n6883), .A2(\mem[240][14] ), .B1(n6174), .B2(
        \mem[246][14] ), .ZN(n4882) );
  AOI22D0 U1103 ( .A1(n6968), .A2(\mem[233][14] ), .B1(n6956), .B2(
        \mem[232][14] ), .ZN(n4880) );
  ND4D0 U1104 ( .A1(n4883), .A2(n4882), .A3(n4881), .A4(n4880), .ZN(n4889) );
  AOI22D0 U1105 ( .A1(n6829), .A2(\mem[230][14] ), .B1(n6639), .B2(
        \mem[231][14] ), .ZN(n4887) );
  AOI22D0 U1106 ( .A1(n6980), .A2(\mem[253][14] ), .B1(n6791), .B2(
        \mem[224][14] ), .ZN(n4886) );
  AOI22D0 U1107 ( .A1(n6991), .A2(\mem[212][14] ), .B1(n6842), .B2(
        \mem[218][14] ), .ZN(n4885) );
  AOI22D0 U1108 ( .A1(n6904), .A2(\mem[211][14] ), .B1(n6760), .B2(
        \mem[237][14] ), .ZN(n4884) );
  ND4D0 U1109 ( .A1(n4887), .A2(n4886), .A3(n4885), .A4(n4884), .ZN(n4888) );
  NR4D0 U1110 ( .A1(n4891), .A2(n4890), .A3(n4889), .A4(n4888), .ZN(n4913) );
  AOI22D0 U1111 ( .A1(n6933), .A2(\mem[225][14] ), .B1(n6836), .B2(
        \mem[202][14] ), .ZN(n4895) );
  AOI22D0 U1112 ( .A1(n6879), .A2(\mem[250][14] ), .B1(n5966), .B2(
        \mem[223][14] ), .ZN(n4894) );
  AOI22D0 U1113 ( .A1(n6759), .A2(\mem[206][14] ), .B1(n6978), .B2(
        \mem[200][14] ), .ZN(n4893) );
  AOI22D0 U1114 ( .A1(n6803), .A2(\mem[247][14] ), .B1(n6707), .B2(
        \mem[215][14] ), .ZN(n4892) );
  ND4D0 U1115 ( .A1(n4895), .A2(n4894), .A3(n4893), .A4(n4892), .ZN(n4911) );
  AOI22D0 U1116 ( .A1(n6790), .A2(\mem[219][14] ), .B1(n6774), .B2(
        \mem[241][14] ), .ZN(n4899) );
  AOI22D0 U1117 ( .A1(n6955), .A2(\mem[213][14] ), .B1(n6871), .B2(
        \mem[249][14] ), .ZN(n4898) );
  AOI22D0 U1118 ( .A1(n6905), .A2(\mem[251][14] ), .B1(n6901), .B2(
        \mem[201][14] ), .ZN(n4897) );
  AOI22D0 U1119 ( .A1(n6892), .A2(\mem[236][14] ), .B1(n6874), .B2(
        \mem[234][14] ), .ZN(n4896) );
  ND4D0 U1120 ( .A1(n4899), .A2(n4898), .A3(n4897), .A4(n4896), .ZN(n4910) );
  AOI22D0 U1121 ( .A1(n6870), .A2(\mem[252][14] ), .B1(n6965), .B2(
        \mem[205][14] ), .ZN(n4903) );
  AOI22D0 U1122 ( .A1(n6525), .A2(\mem[227][14] ), .B1(n6847), .B2(
        \mem[217][14] ), .ZN(n4901) );
  AOI22D0 U1123 ( .A1(n6837), .A2(\mem[207][14] ), .B1(n6828), .B2(
        \mem[248][14] ), .ZN(n4900) );
  ND4D0 U1124 ( .A1(n4903), .A2(n4902), .A3(n4901), .A4(n4900), .ZN(n4909) );
  AOI22D0 U1125 ( .A1(n6802), .A2(\mem[216][14] ), .B1(n6928), .B2(
        \mem[199][14] ), .ZN(n4907) );
  AOI22D0 U1126 ( .A1(n6989), .A2(\mem[198][14] ), .B1(n6754), .B2(
        \mem[197][14] ), .ZN(n4906) );
  AOI22D0 U1127 ( .A1(n6728), .A2(\mem[244][14] ), .B1(n6906), .B2(
        \mem[204][14] ), .ZN(n4905) );
  AOI22D0 U1128 ( .A1(n6890), .A2(\mem[228][14] ), .B1(n6922), .B2(
        \mem[221][14] ), .ZN(n4904) );
  ND4D0 U1129 ( .A1(n4907), .A2(n4906), .A3(n4905), .A4(n4904), .ZN(n4908) );
  NR4D0 U1130 ( .A1(n4911), .A2(n4910), .A3(n4909), .A4(n4908), .ZN(n4912) );
  AOI21D0 U1131 ( .A1(n4913), .A2(n4912), .B(n6945), .ZN(n4957) );
  AOI22D0 U1132 ( .A1(n6861), .A2(\mem[4][14] ), .B1(n6913), .B2(\mem[27][14] ), .ZN(n4917) );
  AOI22D0 U1133 ( .A1(n6928), .A2(\mem[7][14] ), .B1(n6829), .B2(\mem[38][14] ), .ZN(n4916) );
  AOI22D0 U1134 ( .A1(n6880), .A2(\mem[11][14] ), .B1(n6964), .B2(
        \mem[30][14] ), .ZN(n4915) );
  AOI22D0 U1135 ( .A1(n6872), .A2(\mem[6][14] ), .B1(n6916), .B2(\mem[21][14] ), .ZN(n4914) );
  ND4D0 U1136 ( .A1(n4917), .A2(n4916), .A3(n4915), .A4(n4914), .ZN(n4933) );
  AOI22D0 U1137 ( .A1(n6901), .A2(\mem[9][14] ), .B1(n6882), .B2(\mem[15][14] ), .ZN(n4921) );
  AOI22D0 U1138 ( .A1(n6933), .A2(\mem[33][14] ), .B1(n6789), .B2(
        \mem[62][14] ), .ZN(n4920) );
  AOI22D0 U1139 ( .A1(n6952), .A2(\mem[22][14] ), .B1(n6988), .B2(
        \mem[63][14] ), .ZN(n4919) );
  AOI22D0 U1140 ( .A1(n6754), .A2(\mem[5][14] ), .B1(n6738), .B2(\mem[37][14] ), .ZN(n4918) );
  AOI22D0 U1141 ( .A1(n6868), .A2(\mem[43][14] ), .B1(n6863), .B2(
        \mem[55][14] ), .ZN(n4924) );
  AOI22D0 U1142 ( .A1(n6296), .A2(\mem[29][14] ), .B1(n6774), .B2(
        \mem[49][14] ), .ZN(n4923) );
  AOI22D0 U1143 ( .A1(n6860), .A2(\mem[35][14] ), .B1(n6904), .B2(
        \mem[19][14] ), .ZN(n4922) );
  ND4D0 U1144 ( .A1(n4925), .A2(n4924), .A3(n4923), .A4(n4922), .ZN(n4931) );
  AOI22D0 U1145 ( .A1(n6980), .A2(\mem[61][14] ), .B1(n6926), .B2(\mem[1][14] ), .ZN(n4929) );
  AOI22D0 U1146 ( .A1(n6917), .A2(\mem[46][14] ), .B1(n6991), .B2(
        \mem[20][14] ), .ZN(n4928) );
  AOI22D0 U1147 ( .A1(n6448), .A2(\mem[0][14] ), .B1(n6978), .B2(\mem[8][14] ), 
        .ZN(n4927) );
  AOI22D0 U1148 ( .A1(n6759), .A2(\mem[14][14] ), .B1(n6760), .B2(
        \mem[45][14] ), .ZN(n4926) );
  ND4D0 U1149 ( .A1(n4929), .A2(n4928), .A3(n4927), .A4(n4926), .ZN(n4930) );
  NR4D0 U1150 ( .A1(n4933), .A2(n4932), .A3(n4931), .A4(n4930), .ZN(n4955) );
  AOI22D0 U1151 ( .A1(n6883), .A2(\mem[48][14] ), .B1(n6970), .B2(
        \mem[16][14] ), .ZN(n4937) );
  AOI22D0 U1152 ( .A1(n6784), .A2(\mem[28][14] ), .B1(n6639), .B2(
        \mem[39][14] ), .ZN(n4936) );
  AOI22D0 U1153 ( .A1(n6924), .A2(\mem[32][14] ), .B1(n6707), .B2(
        \mem[23][14] ), .ZN(n4935) );
  AOI22D0 U1154 ( .A1(n6680), .A2(\mem[31][14] ), .B1(n6847), .B2(
        \mem[25][14] ), .ZN(n4934) );
  ND4D0 U1155 ( .A1(n4937), .A2(n4936), .A3(n4935), .A4(n4934), .ZN(n4953) );
  AOI22D0 U1156 ( .A1(n6993), .A2(\mem[53][14] ), .B1(n6957), .B2(
        \mem[57][14] ), .ZN(n4941) );
  AOI22D0 U1157 ( .A1(n6870), .A2(\mem[60][14] ), .B1(n6874), .B2(
        \mem[42][14] ), .ZN(n4940) );
  AOI22D0 U1158 ( .A1(n6891), .A2(\mem[26][14] ), .B1(n6936), .B2(
        \mem[17][14] ), .ZN(n4939) );
  ND4D0 U1159 ( .A1(n4941), .A2(n4940), .A3(n4939), .A4(n4938), .ZN(n4952) );
  AOI22D0 U1160 ( .A1(n6959), .A2(\mem[3][14] ), .B1(n6992), .B2(\mem[54][14] ), .ZN(n4945) );
  AOI22D0 U1161 ( .A1(n6890), .A2(\mem[36][14] ), .B1(n6491), .B2(
        \mem[51][14] ), .ZN(n4944) );
  AOI22D0 U1162 ( .A1(n6905), .A2(\mem[59][14] ), .B1(n6542), .B2(
        \mem[18][14] ), .ZN(n4943) );
  AOI22D0 U1163 ( .A1(n6179), .A2(\mem[47][14] ), .B1(n6698), .B2(\mem[2][14] ), .ZN(n4942) );
  ND4D0 U1164 ( .A1(n4945), .A2(n4944), .A3(n4943), .A4(n4942), .ZN(n4951) );
  AOI22D0 U1165 ( .A1(n6912), .A2(\mem[56][14] ), .B1(n6906), .B2(
        \mem[12][14] ), .ZN(n4949) );
  AOI22D0 U1166 ( .A1(n6934), .A2(\mem[24][14] ), .B1(n6956), .B2(
        \mem[40][14] ), .ZN(n4948) );
  AOI22D0 U1167 ( .A1(n6892), .A2(\mem[44][14] ), .B1(n6879), .B2(
        \mem[58][14] ), .ZN(n4947) );
  AOI22D0 U1168 ( .A1(n6923), .A2(\mem[34][14] ), .B1(n6836), .B2(
        \mem[10][14] ), .ZN(n4946) );
  ND4D0 U1169 ( .A1(n4949), .A2(n4948), .A3(n4947), .A4(n4946), .ZN(n4950) );
  NR4D0 U1170 ( .A1(n4953), .A2(n4952), .A3(n4951), .A4(n4950), .ZN(n4954) );
  AOI211D0 U1171 ( .A1(n6951), .A2(n4958), .B(n4957), .C(n4956), .ZN(n4980) );
  AOI22D0 U1172 ( .A1(n6928), .A2(\mem[71][14] ), .B1(n6923), .B2(
        \mem[98][14] ), .ZN(n4962) );
  AOI22D0 U1173 ( .A1(n6907), .A2(\mem[67][14] ), .B1(n6835), .B2(
        \mem[68][14] ), .ZN(n4961) );
  AOI22D0 U1174 ( .A1(n6680), .A2(\mem[95][14] ), .B1(n6491), .B2(
        \mem[115][14] ), .ZN(n4959) );
  ND4D0 U1175 ( .A1(n4962), .A2(n4961), .A3(n4960), .A4(n4959), .ZN(n4978) );
  AOI22D0 U1176 ( .A1(n6814), .A2(\mem[65][14] ), .B1(n6847), .B2(
        \mem[89][14] ), .ZN(n4966) );
  AOI22D0 U1177 ( .A1(n6784), .A2(\mem[92][14] ), .B1(n6965), .B2(
        \mem[77][14] ), .ZN(n4965) );
  AOI22D0 U1178 ( .A1(n6733), .A2(\mem[122][14] ), .B1(n6828), .B2(
        \mem[120][14] ), .ZN(n4964) );
  AOI22D0 U1179 ( .A1(n6953), .A2(\mem[111][14] ), .B1(n6891), .B2(
        \mem[90][14] ), .ZN(n4963) );
  ND4D0 U1180 ( .A1(n4966), .A2(n4965), .A3(n4964), .A4(n4963), .ZN(n4977) );
  AOI22D0 U1181 ( .A1(n6990), .A2(\mem[76][14] ), .B1(n6774), .B2(
        \mem[113][14] ), .ZN(n4970) );
  AOI22D0 U1182 ( .A1(n6995), .A2(\mem[87][14] ), .B1(n6738), .B2(
        \mem[101][14] ), .ZN(n4969) );
  AOI22D0 U1183 ( .A1(n6969), .A2(\mem[82][14] ), .B1(n6658), .B2(
        \mem[114][14] ), .ZN(n4968) );
  AOI22D0 U1184 ( .A1(n6971), .A2(\mem[102][14] ), .B1(n6748), .B2(
        \mem[105][14] ), .ZN(n4967) );
  ND4D0 U1185 ( .A1(n4970), .A2(n4969), .A3(n4968), .A4(n4967), .ZN(n4976) );
  AOI22D0 U1186 ( .A1(n6802), .A2(\mem[88][14] ), .B1(n6933), .B2(
        \mem[97][14] ), .ZN(n4974) );
  AOI22D0 U1187 ( .A1(n6913), .A2(\mem[91][14] ), .B1(n6936), .B2(
        \mem[81][14] ), .ZN(n4973) );
  AOI22D0 U1188 ( .A1(n6868), .A2(\mem[107][14] ), .B1(n6698), .B2(
        \mem[66][14] ), .ZN(n4972) );
  AOI22D0 U1189 ( .A1(n6881), .A2(\mem[80][14] ), .B1(n6789), .B2(
        \mem[126][14] ), .ZN(n4971) );
  ND4D0 U1190 ( .A1(n4974), .A2(n4973), .A3(n4972), .A4(n4971), .ZN(n4975) );
  NR4D0 U1191 ( .A1(n4978), .A2(n4977), .A3(n4976), .A4(n4975), .ZN(n4979) );
  AOI32D0 U1192 ( .A1(n4981), .A2(n4980), .A3(n4979), .B1(n7004), .B2(n4980), 
        .ZN(dout[14]) );
  AOI22D0 U1193 ( .A1(n6933), .A2(\mem[33][12] ), .B1(n6847), .B2(
        \mem[25][12] ), .ZN(n4985) );
  AOI22D0 U1194 ( .A1(n6542), .A2(\mem[18][12] ), .B1(n6881), .B2(
        \mem[16][12] ), .ZN(n4984) );
  AOI22D0 U1195 ( .A1(n6829), .A2(\mem[38][12] ), .B1(n6639), .B2(
        \mem[39][12] ), .ZN(n4983) );
  AOI22D0 U1196 ( .A1(n6870), .A2(\mem[60][12] ), .B1(n6774), .B2(
        \mem[49][12] ), .ZN(n4982) );
  ND4D0 U1197 ( .A1(n4985), .A2(n4984), .A3(n4983), .A4(n4982), .ZN(n5001) );
  AOI22D0 U1198 ( .A1(n6880), .A2(\mem[11][12] ), .B1(n6904), .B2(
        \mem[19][12] ), .ZN(n4989) );
  AOI22D0 U1199 ( .A1(n6803), .A2(\mem[55][12] ), .B1(n6982), .B2(\mem[2][12] ), .ZN(n4988) );
  AOI22D0 U1200 ( .A1(n6759), .A2(\mem[14][12] ), .B1(n6491), .B2(
        \mem[51][12] ), .ZN(n4987) );
  ND4D0 U1201 ( .A1(n4989), .A2(n4988), .A3(n4987), .A4(n4986), .ZN(n5000) );
  AOI22D0 U1202 ( .A1(n6784), .A2(\mem[28][12] ), .B1(n6913), .B2(
        \mem[27][12] ), .ZN(n4993) );
  AOI22D0 U1203 ( .A1(n6955), .A2(\mem[21][12] ), .B1(n6992), .B2(
        \mem[54][12] ), .ZN(n4992) );
  AOI22D0 U1204 ( .A1(n6872), .A2(\mem[6][12] ), .B1(n6874), .B2(\mem[42][12] ), .ZN(n4991) );
  AOI22D0 U1205 ( .A1(n6680), .A2(\mem[31][12] ), .B1(n6936), .B2(
        \mem[17][12] ), .ZN(n4990) );
  ND4D0 U1206 ( .A1(n4993), .A2(n4992), .A3(n4991), .A4(n4990), .ZN(n4999) );
  AOI22D0 U1207 ( .A1(n6871), .A2(\mem[57][12] ), .B1(n6964), .B2(
        \mem[30][12] ), .ZN(n4997) );
  AOI22D0 U1208 ( .A1(n6747), .A2(\mem[20][12] ), .B1(n6922), .B2(
        \mem[29][12] ), .ZN(n4996) );
  AOI22D0 U1209 ( .A1(n6928), .A2(\mem[7][12] ), .B1(n6860), .B2(\mem[35][12] ), .ZN(n4995) );
  AOI22D0 U1210 ( .A1(n6995), .A2(\mem[23][12] ), .B1(n6748), .B2(
        \mem[41][12] ), .ZN(n4994) );
  ND4D0 U1211 ( .A1(n4997), .A2(n4996), .A3(n4995), .A4(n4994), .ZN(n4998) );
  NR4D0 U1212 ( .A1(n5001), .A2(n5000), .A3(n4999), .A4(n4998), .ZN(n5153) );
  AOI22D0 U1213 ( .A1(n6967), .A2(\mem[167][12] ), .B1(n6828), .B2(
        \mem[184][12] ), .ZN(n5005) );
  AOI22D0 U1214 ( .A1(n6952), .A2(\mem[150][12] ), .B1(n6901), .B2(
        \mem[137][12] ), .ZN(n5004) );
  AOI22D0 U1215 ( .A1(n6814), .A2(\mem[129][12] ), .B1(n6882), .B2(
        \mem[143][12] ), .ZN(n5003) );
  AOI22D0 U1216 ( .A1(n6966), .A2(\mem[178][12] ), .B1(n6964), .B2(
        \mem[158][12] ), .ZN(n5002) );
  ND4D0 U1217 ( .A1(n5005), .A2(n5004), .A3(n5003), .A4(n5002), .ZN(n5021) );
  AOI22D0 U1218 ( .A1(n6890), .A2(\mem[164][12] ), .B1(n6983), .B2(
        \mem[176][12] ), .ZN(n5009) );
  AOI22D0 U1219 ( .A1(n6448), .A2(\mem[128][12] ), .B1(n6707), .B2(
        \mem[151][12] ), .ZN(n5008) );
  AOI22D0 U1220 ( .A1(n6922), .A2(\mem[157][12] ), .B1(n6174), .B2(
        \mem[182][12] ), .ZN(n5007) );
  AOI22D0 U1221 ( .A1(n6749), .A2(\mem[171][12] ), .B1(n6842), .B2(
        \mem[154][12] ), .ZN(n5006) );
  ND4D0 U1222 ( .A1(n5009), .A2(n5008), .A3(n5007), .A4(n5006), .ZN(n5020) );
  AOI22D0 U1223 ( .A1(n6165), .A2(\mem[174][12] ), .B1(n6804), .B2(
        \mem[147][12] ), .ZN(n5013) );
  AOI22D0 U1224 ( .A1(n6530), .A2(\mem[187][12] ), .B1(n6988), .B2(
        \mem[191][12] ), .ZN(n5012) );
  AOI22D0 U1225 ( .A1(n6953), .A2(\mem[175][12] ), .B1(n6863), .B2(
        \mem[183][12] ), .ZN(n5011) );
  AOI22D0 U1226 ( .A1(n6925), .A2(\mem[173][12] ), .B1(n6738), .B2(
        \mem[165][12] ), .ZN(n5010) );
  ND4D0 U1227 ( .A1(n5013), .A2(n5012), .A3(n5011), .A4(n5010), .ZN(n5019) );
  AOI22D0 U1228 ( .A1(n6802), .A2(\mem[152][12] ), .B1(n6994), .B2(
        \mem[190][12] ), .ZN(n5017) );
  AOI22D0 U1229 ( .A1(n6847), .A2(\mem[153][12] ), .B1(n6748), .B2(
        \mem[169][12] ), .ZN(n5016) );
  AOI22D0 U1230 ( .A1(n6959), .A2(\mem[131][12] ), .B1(n6860), .B2(
        \mem[163][12] ), .ZN(n5014) );
  ND4D0 U1231 ( .A1(n5017), .A2(n5016), .A3(n5015), .A4(n5014), .ZN(n5018) );
  NR4D0 U1232 ( .A1(n5021), .A2(n5020), .A3(n5019), .A4(n5018), .ZN(n5043) );
  AOI22D0 U1233 ( .A1(n6977), .A2(\mem[161][12] ), .B1(n6906), .B2(
        \mem[140][12] ), .ZN(n5025) );
  AOI22D0 U1234 ( .A1(n6981), .A2(\mem[188][12] ), .B1(n6991), .B2(
        \mem[148][12] ), .ZN(n5024) );
  AOI22D0 U1235 ( .A1(n6680), .A2(\mem[159][12] ), .B1(n6728), .B2(
        \mem[180][12] ), .ZN(n5023) );
  AOI22D0 U1236 ( .A1(n6784), .A2(\mem[156][12] ), .B1(n6969), .B2(
        \mem[146][12] ), .ZN(n5022) );
  ND4D0 U1237 ( .A1(n5025), .A2(n5024), .A3(n5023), .A4(n5022), .ZN(n5041) );
  AOI22D0 U1238 ( .A1(n6759), .A2(\mem[142][12] ), .B1(n6965), .B2(
        \mem[141][12] ), .ZN(n5029) );
  AOI22D0 U1239 ( .A1(n6775), .A2(\mem[172][12] ), .B1(n6774), .B2(
        \mem[177][12] ), .ZN(n5028) );
  AOI22D0 U1240 ( .A1(n6325), .A2(\mem[139][12] ), .B1(n6989), .B2(
        \mem[134][12] ), .ZN(n5027) );
  AOI22D0 U1241 ( .A1(n6754), .A2(\mem[133][12] ), .B1(n6903), .B2(
        \mem[179][12] ), .ZN(n5026) );
  ND4D0 U1242 ( .A1(n5029), .A2(n5028), .A3(n5027), .A4(n5026), .ZN(n5040) );
  AOI22D0 U1243 ( .A1(n6830), .A2(\mem[135][12] ), .B1(n6956), .B2(
        \mem[168][12] ), .ZN(n5033) );
  AOI22D0 U1244 ( .A1(n6835), .A2(\mem[132][12] ), .B1(n6698), .B2(
        \mem[130][12] ), .ZN(n5032) );
  AOI22D0 U1245 ( .A1(n6971), .A2(\mem[166][12] ), .B1(n6791), .B2(
        \mem[160][12] ), .ZN(n5031) );
  AOI22D0 U1246 ( .A1(n6727), .A2(\mem[170][12] ), .B1(n6978), .B2(
        \mem[136][12] ), .ZN(n5030) );
  ND4D0 U1247 ( .A1(n5033), .A2(n5032), .A3(n5031), .A4(n5030), .ZN(n5039) );
  AOI22D0 U1248 ( .A1(n6955), .A2(\mem[149][12] ), .B1(n6936), .B2(
        \mem[145][12] ), .ZN(n5037) );
  AOI22D0 U1249 ( .A1(n6879), .A2(\mem[186][12] ), .B1(n6957), .B2(
        \mem[185][12] ), .ZN(n5035) );
  AOI22D0 U1250 ( .A1(n6980), .A2(\mem[189][12] ), .B1(n6954), .B2(
        \mem[138][12] ), .ZN(n5034) );
  ND4D0 U1251 ( .A1(n5037), .A2(n5036), .A3(n5035), .A4(n5034), .ZN(n5038) );
  NR4D0 U1252 ( .A1(n5041), .A2(n5040), .A3(n5039), .A4(n5038), .ZN(n5042) );
  AOI22D0 U1253 ( .A1(n6917), .A2(\mem[110][12] ), .B1(n6936), .B2(
        \mem[81][12] ), .ZN(n5047) );
  AOI22D0 U1254 ( .A1(n6969), .A2(\mem[82][12] ), .B1(n6863), .B2(
        \mem[119][12] ), .ZN(n5046) );
  AOI22D0 U1255 ( .A1(n6977), .A2(\mem[97][12] ), .B1(n6874), .B2(
        \mem[106][12] ), .ZN(n5045) );
  AOI22D0 U1256 ( .A1(n6881), .A2(\mem[80][12] ), .B1(n6748), .B2(
        \mem[105][12] ), .ZN(n5044) );
  ND4D0 U1257 ( .A1(n5047), .A2(n5046), .A3(n5045), .A4(n5044), .ZN(n5063) );
  AOI22D0 U1258 ( .A1(n6747), .A2(\mem[84][12] ), .B1(n6978), .B2(
        \mem[72][12] ), .ZN(n5051) );
  AOI22D0 U1259 ( .A1(n6784), .A2(\mem[92][12] ), .B1(n6906), .B2(
        \mem[76][12] ), .ZN(n5050) );
  AOI22D0 U1260 ( .A1(n6922), .A2(\mem[93][12] ), .B1(n6955), .B2(
        \mem[85][12] ), .ZN(n5049) );
  AOI22D0 U1261 ( .A1(n6819), .A2(\mem[125][12] ), .B1(n6924), .B2(
        \mem[96][12] ), .ZN(n5048) );
  ND4D0 U1262 ( .A1(n5051), .A2(n5050), .A3(n5049), .A4(n5048), .ZN(n5062) );
  AOI22D0 U1263 ( .A1(n6530), .A2(\mem[123][12] ), .B1(n6847), .B2(
        \mem[89][12] ), .ZN(n5055) );
  AOI22D0 U1264 ( .A1(n6868), .A2(\mem[107][12] ), .B1(n6880), .B2(
        \mem[75][12] ), .ZN(n5054) );
  AOI22D0 U1265 ( .A1(n6890), .A2(\mem[100][12] ), .B1(n6971), .B2(
        \mem[102][12] ), .ZN(n5053) );
  AOI22D0 U1266 ( .A1(n6448), .A2(\mem[64][12] ), .B1(n6993), .B2(
        \mem[117][12] ), .ZN(n5052) );
  ND4D0 U1267 ( .A1(n5055), .A2(n5054), .A3(n5053), .A4(n5052), .ZN(n5061) );
  AOI22D0 U1268 ( .A1(n6981), .A2(\mem[124][12] ), .B1(n6979), .B2(
        \mem[78][12] ), .ZN(n5058) );
  AOI22D0 U1269 ( .A1(n6775), .A2(\mem[108][12] ), .B1(n6879), .B2(
        \mem[122][12] ), .ZN(n5057) );
  AOI22D0 U1270 ( .A1(n6994), .A2(\mem[126][12] ), .B1(n6774), .B2(
        \mem[113][12] ), .ZN(n5056) );
  ND4D0 U1271 ( .A1(n5059), .A2(n5058), .A3(n5057), .A4(n5056), .ZN(n5060) );
  NR4D0 U1272 ( .A1(n5063), .A2(n5062), .A3(n5061), .A4(n5060), .ZN(n5085) );
  AOI22D0 U1273 ( .A1(n6907), .A2(\mem[67][12] ), .B1(n6836), .B2(
        \mem[74][12] ), .ZN(n5067) );
  AOI22D0 U1274 ( .A1(n6809), .A2(\mem[73][12] ), .B1(n6828), .B2(
        \mem[120][12] ), .ZN(n5066) );
  AOI22D0 U1275 ( .A1(n6790), .A2(\mem[91][12] ), .B1(n6982), .B2(
        \mem[66][12] ), .ZN(n5065) );
  AOI22D0 U1276 ( .A1(n6680), .A2(\mem[95][12] ), .B1(n6965), .B2(
        \mem[77][12] ), .ZN(n5064) );
  ND4D0 U1277 ( .A1(n5067), .A2(n5066), .A3(n5065), .A4(n5064), .ZN(n5083) );
  AOI22D0 U1278 ( .A1(n6923), .A2(\mem[98][12] ), .B1(n6988), .B2(
        \mem[127][12] ), .ZN(n5071) );
  AOI22D0 U1279 ( .A1(n6525), .A2(\mem[99][12] ), .B1(n6871), .B2(
        \mem[121][12] ), .ZN(n5070) );
  AOI22D0 U1280 ( .A1(n6658), .A2(\mem[114][12] ), .B1(n6904), .B2(
        \mem[83][12] ), .ZN(n5069) );
  AOI22D0 U1281 ( .A1(n6903), .A2(\mem[115][12] ), .B1(n6964), .B2(
        \mem[94][12] ), .ZN(n5068) );
  ND4D0 U1282 ( .A1(n5071), .A2(n5070), .A3(n5069), .A4(n5068), .ZN(n5082) );
  AOI22D0 U1283 ( .A1(n6883), .A2(\mem[112][12] ), .B1(n6728), .B2(
        \mem[116][12] ), .ZN(n5075) );
  AOI22D0 U1284 ( .A1(n6814), .A2(\mem[65][12] ), .B1(n6835), .B2(
        \mem[68][12] ), .ZN(n5074) );
  AOI22D0 U1285 ( .A1(n6967), .A2(\mem[103][12] ), .B1(n6992), .B2(
        \mem[118][12] ), .ZN(n5073) );
  AOI22D0 U1286 ( .A1(n6952), .A2(\mem[86][12] ), .B1(n6882), .B2(
        \mem[79][12] ), .ZN(n5079) );
  AOI22D0 U1287 ( .A1(n6995), .A2(\mem[87][12] ), .B1(n6956), .B2(
        \mem[104][12] ), .ZN(n5078) );
  AOI22D0 U1288 ( .A1(n6934), .A2(\mem[88][12] ), .B1(n6738), .B2(
        \mem[101][12] ), .ZN(n5077) );
  AOI22D0 U1289 ( .A1(n6872), .A2(\mem[70][12] ), .B1(n6754), .B2(
        \mem[69][12] ), .ZN(n5076) );
  ND4D0 U1290 ( .A1(n5079), .A2(n5078), .A3(n5077), .A4(n5076), .ZN(n5080) );
  NR4D0 U1291 ( .A1(n5083), .A2(n5082), .A3(n5081), .A4(n5080), .ZN(n5084) );
  AOI21D0 U1292 ( .A1(n5085), .A2(n5084), .B(n7004), .ZN(n5129) );
  AOI22D0 U1293 ( .A1(n6830), .A2(\mem[199][12] ), .B1(n6978), .B2(
        \mem[200][12] ), .ZN(n5089) );
  AOI22D0 U1294 ( .A1(n6861), .A2(\mem[196][12] ), .B1(n6922), .B2(
        \mem[221][12] ), .ZN(n5088) );
  AOI22D0 U1295 ( .A1(n6784), .A2(\mem[220][12] ), .B1(n6956), .B2(
        \mem[232][12] ), .ZN(n5087) );
  AOI22D0 U1296 ( .A1(n6868), .A2(\mem[235][12] ), .B1(n6760), .B2(
        \mem[237][12] ), .ZN(n5086) );
  ND4D0 U1297 ( .A1(n5089), .A2(n5088), .A3(n5087), .A4(n5086), .ZN(n5105) );
  AOI22D0 U1298 ( .A1(n6958), .A2(\mem[209][12] ), .B1(n6836), .B2(
        \mem[202][12] ), .ZN(n5093) );
  AOI22D0 U1299 ( .A1(n6903), .A2(\mem[243][12] ), .B1(n6791), .B2(
        \mem[224][12] ), .ZN(n5092) );
  AOI22D0 U1300 ( .A1(n6542), .A2(\mem[210][12] ), .B1(n6863), .B2(
        \mem[247][12] ), .ZN(n5091) );
  AOI22D0 U1301 ( .A1(n6993), .A2(\mem[245][12] ), .B1(n6992), .B2(
        \mem[246][12] ), .ZN(n5090) );
  ND4D0 U1302 ( .A1(n5093), .A2(n5092), .A3(n5091), .A4(n5090), .ZN(n5104) );
  AOI22D0 U1303 ( .A1(n5966), .A2(\mem[223][12] ), .B1(n6789), .B2(
        \mem[254][12] ), .ZN(n5097) );
  AOI22D0 U1304 ( .A1(n6879), .A2(\mem[250][12] ), .B1(n6966), .B2(
        \mem[242][12] ), .ZN(n5096) );
  AOI22D0 U1305 ( .A1(n6917), .A2(\mem[238][12] ), .B1(n6959), .B2(
        \mem[195][12] ), .ZN(n5094) );
  ND4D0 U1306 ( .A1(n5097), .A2(n5096), .A3(n5095), .A4(n5094), .ZN(n5103) );
  AOI22D0 U1307 ( .A1(n6880), .A2(\mem[203][12] ), .B1(n6957), .B2(
        \mem[249][12] ), .ZN(n5101) );
  AOI22D0 U1308 ( .A1(n6952), .A2(\mem[214][12] ), .B1(n6698), .B2(
        \mem[194][12] ), .ZN(n5100) );
  AOI22D0 U1309 ( .A1(n6819), .A2(\mem[253][12] ), .B1(n6804), .B2(
        \mem[211][12] ), .ZN(n5099) );
  AOI22D0 U1310 ( .A1(n6882), .A2(\mem[207][12] ), .B1(n6964), .B2(
        \mem[222][12] ), .ZN(n5098) );
  ND4D0 U1311 ( .A1(n5101), .A2(n5100), .A3(n5099), .A4(n5098), .ZN(n5102) );
  NR4D0 U1312 ( .A1(n5105), .A2(n5104), .A3(n5103), .A4(n5102), .ZN(n5127) );
  AOI22D0 U1313 ( .A1(n6530), .A2(\mem[251][12] ), .B1(n6933), .B2(
        \mem[225][12] ), .ZN(n5109) );
  AOI22D0 U1314 ( .A1(n6448), .A2(\mem[192][12] ), .B1(n6842), .B2(
        \mem[218][12] ), .ZN(n5108) );
  AOI22D0 U1315 ( .A1(n6747), .A2(\mem[212][12] ), .B1(n6869), .B2(
        \mem[241][12] ), .ZN(n5107) );
  AOI22D0 U1316 ( .A1(n6870), .A2(\mem[252][12] ), .B1(n6983), .B2(
        \mem[240][12] ), .ZN(n5106) );
  ND4D0 U1317 ( .A1(n5109), .A2(n5108), .A3(n5107), .A4(n5106), .ZN(n5125) );
  AOI22D0 U1318 ( .A1(n6814), .A2(\mem[193][12] ), .B1(n6923), .B2(
        \mem[226][12] ), .ZN(n5113) );
  AOI22D0 U1319 ( .A1(n6914), .A2(\mem[197][12] ), .B1(n6965), .B2(
        \mem[205][12] ), .ZN(n5112) );
  AOI22D0 U1320 ( .A1(n6775), .A2(\mem[236][12] ), .B1(n6639), .B2(
        \mem[231][12] ), .ZN(n5111) );
  AOI22D0 U1321 ( .A1(n6913), .A2(\mem[219][12] ), .B1(n6902), .B2(
        \mem[229][12] ), .ZN(n5110) );
  ND4D0 U1322 ( .A1(n5113), .A2(n5112), .A3(n5111), .A4(n5110), .ZN(n5124) );
  AOI22D0 U1323 ( .A1(n6970), .A2(\mem[208][12] ), .B1(n6906), .B2(
        \mem[204][12] ), .ZN(n5117) );
  AOI22D0 U1324 ( .A1(n6727), .A2(\mem[234][12] ), .B1(n6968), .B2(
        \mem[233][12] ), .ZN(n5115) );
  AOI22D0 U1325 ( .A1(n6995), .A2(\mem[215][12] ), .B1(n6728), .B2(
        \mem[244][12] ), .ZN(n5114) );
  ND4D0 U1326 ( .A1(n5117), .A2(n5116), .A3(n5115), .A4(n5114), .ZN(n5123) );
  AOI22D0 U1327 ( .A1(n6802), .A2(\mem[216][12] ), .B1(n6828), .B2(
        \mem[248][12] ), .ZN(n5121) );
  AOI22D0 U1328 ( .A1(n6525), .A2(\mem[227][12] ), .B1(n6971), .B2(
        \mem[230][12] ), .ZN(n5120) );
  AOI22D0 U1329 ( .A1(n6890), .A2(\mem[228][12] ), .B1(n6989), .B2(
        \mem[198][12] ), .ZN(n5119) );
  AOI22D0 U1330 ( .A1(n6847), .A2(\mem[217][12] ), .B1(n6916), .B2(
        \mem[213][12] ), .ZN(n5118) );
  ND4D0 U1331 ( .A1(n5121), .A2(n5120), .A3(n5119), .A4(n5118), .ZN(n5122) );
  NR4D0 U1332 ( .A1(n5125), .A2(n5124), .A3(n5123), .A4(n5122), .ZN(n5126) );
  AOI21D0 U1333 ( .A1(n5127), .A2(n5126), .B(n6945), .ZN(n5128) );
  AOI211D0 U1334 ( .A1(n6951), .A2(n5130), .B(n5129), .C(n5128), .ZN(n5152) );
  AOI22D0 U1335 ( .A1(n6835), .A2(\mem[4][12] ), .B1(n6993), .B2(\mem[53][12] ), .ZN(n5133) );
  AOI22D0 U1336 ( .A1(n6923), .A2(\mem[34][12] ), .B1(n6760), .B2(
        \mem[45][12] ), .ZN(n5132) );
  AOI22D0 U1337 ( .A1(n6980), .A2(\mem[61][12] ), .B1(n6892), .B2(
        \mem[44][12] ), .ZN(n5131) );
  ND4D0 U1338 ( .A1(n5134), .A2(n5133), .A3(n5132), .A4(n5131), .ZN(n5150) );
  AOI22D0 U1339 ( .A1(n6907), .A2(\mem[3][12] ), .B1(n6924), .B2(\mem[32][12] ), .ZN(n5138) );
  AOI22D0 U1340 ( .A1(n6953), .A2(\mem[47][12] ), .B1(n6836), .B2(
        \mem[10][12] ), .ZN(n5137) );
  AOI22D0 U1341 ( .A1(n6915), .A2(\mem[13][12] ), .B1(n6978), .B2(\mem[8][12] ), .ZN(n5136) );
  AOI22D0 U1342 ( .A1(n6814), .A2(\mem[1][12] ), .B1(n6988), .B2(\mem[63][12] ), .ZN(n5135) );
  ND4D0 U1343 ( .A1(n5138), .A2(n5137), .A3(n5136), .A4(n5135), .ZN(n5149) );
  AOI22D0 U1344 ( .A1(n6802), .A2(\mem[24][12] ), .B1(n6809), .B2(\mem[9][12] ), .ZN(n5142) );
  AOI22D0 U1345 ( .A1(n6773), .A2(\mem[36][12] ), .B1(n6990), .B2(
        \mem[12][12] ), .ZN(n5141) );
  AOI22D0 U1346 ( .A1(n6448), .A2(\mem[0][12] ), .B1(n6842), .B2(\mem[26][12] ), .ZN(n5140) );
  AOI22D0 U1347 ( .A1(n6879), .A2(\mem[58][12] ), .B1(n6828), .B2(
        \mem[56][12] ), .ZN(n5139) );
  ND4D0 U1348 ( .A1(n5142), .A2(n5141), .A3(n5140), .A4(n5139), .ZN(n5148) );
  AOI22D0 U1349 ( .A1(n6868), .A2(\mem[43][12] ), .B1(n6862), .B2(
        \mem[40][12] ), .ZN(n5146) );
  AOI22D0 U1350 ( .A1(n6952), .A2(\mem[22][12] ), .B1(n6983), .B2(
        \mem[48][12] ), .ZN(n5145) );
  AOI22D0 U1351 ( .A1(n6914), .A2(\mem[5][12] ), .B1(n6738), .B2(\mem[37][12] ), .ZN(n5144) );
  ND4D0 U1352 ( .A1(n5146), .A2(n5145), .A3(n5144), .A4(n5143), .ZN(n5147) );
  NR4D0 U1353 ( .A1(n5150), .A2(n5149), .A3(n5148), .A4(n5147), .ZN(n5151) );
  AOI32D0 U1354 ( .A1(n5153), .A2(n5152), .A3(n5151), .B1(n6856), .B2(n5152), 
        .ZN(dout[12]) );
  AOI22D0 U1355 ( .A1(n6759), .A2(\mem[14][11] ), .B1(n6912), .B2(
        \mem[56][11] ), .ZN(n5157) );
  AOI22D0 U1356 ( .A1(n6922), .A2(\mem[29][11] ), .B1(n6789), .B2(
        \mem[62][11] ), .ZN(n5156) );
  AOI22D0 U1357 ( .A1(n6933), .A2(\mem[33][11] ), .B1(n6842), .B2(
        \mem[26][11] ), .ZN(n5155) );
  AOI22D0 U1358 ( .A1(n6907), .A2(\mem[3][11] ), .B1(n6754), .B2(\mem[5][11] ), 
        .ZN(n5154) );
  ND4D0 U1359 ( .A1(n5157), .A2(n5156), .A3(n5155), .A4(n5154), .ZN(n5173) );
  AOI22D0 U1360 ( .A1(n6917), .A2(\mem[46][11] ), .B1(n6991), .B2(
        \mem[20][11] ), .ZN(n5161) );
  AOI22D0 U1361 ( .A1(n6802), .A2(\mem[24][11] ), .B1(n6563), .B2(\mem[8][11] ), .ZN(n5160) );
  AOI22D0 U1362 ( .A1(n6784), .A2(\mem[28][11] ), .B1(n6935), .B2(
        \mem[63][11] ), .ZN(n5159) );
  AOI22D0 U1363 ( .A1(n6803), .A2(\mem[55][11] ), .B1(n6965), .B2(
        \mem[13][11] ), .ZN(n5158) );
  ND4D0 U1364 ( .A1(n5161), .A2(n5160), .A3(n5159), .A4(n5158), .ZN(n5172) );
  AOI22D0 U1365 ( .A1(n6819), .A2(\mem[61][11] ), .B1(n6639), .B2(
        \mem[39][11] ), .ZN(n5165) );
  AOI22D0 U1366 ( .A1(n6970), .A2(\mem[16][11] ), .B1(n6901), .B2(\mem[9][11] ), .ZN(n5164) );
  AOI22D0 U1367 ( .A1(n6871), .A2(\mem[57][11] ), .B1(n6873), .B2(
        \mem[30][11] ), .ZN(n5163) );
  AOI22D0 U1368 ( .A1(n6924), .A2(\mem[32][11] ), .B1(n6992), .B2(
        \mem[54][11] ), .ZN(n5162) );
  ND4D0 U1369 ( .A1(n5165), .A2(n5164), .A3(n5163), .A4(n5162), .ZN(n5171) );
  AOI22D0 U1370 ( .A1(n6525), .A2(\mem[35][11] ), .B1(n6913), .B2(
        \mem[27][11] ), .ZN(n5169) );
  AOI22D0 U1371 ( .A1(n6872), .A2(\mem[6][11] ), .B1(n6888), .B2(\mem[0][11] ), 
        .ZN(n5167) );
  AOI22D0 U1372 ( .A1(n6728), .A2(\mem[52][11] ), .B1(n6902), .B2(
        \mem[37][11] ), .ZN(n5166) );
  ND4D0 U1373 ( .A1(n5169), .A2(n5168), .A3(n5167), .A4(n5166), .ZN(n5170) );
  NR4D0 U1374 ( .A1(n5173), .A2(n5172), .A3(n5171), .A4(n5170), .ZN(n5325) );
  AOI22D0 U1375 ( .A1(n6803), .A2(\mem[183][11] ), .B1(n6738), .B2(
        \mem[165][11] ), .ZN(n5177) );
  AOI22D0 U1376 ( .A1(n6907), .A2(\mem[131][11] ), .B1(n6965), .B2(
        \mem[141][11] ), .ZN(n5176) );
  AOI22D0 U1377 ( .A1(n6881), .A2(\mem[144][11] ), .B1(n6958), .B2(
        \mem[145][11] ), .ZN(n5175) );
  AOI22D0 U1378 ( .A1(n6952), .A2(\mem[150][11] ), .B1(n6991), .B2(
        \mem[148][11] ), .ZN(n5174) );
  ND4D0 U1379 ( .A1(n5177), .A2(n5176), .A3(n5175), .A4(n5174), .ZN(n5193) );
  AOI22D0 U1380 ( .A1(n6814), .A2(\mem[129][11] ), .B1(n6925), .B2(
        \mem[173][11] ), .ZN(n5181) );
  AOI22D0 U1381 ( .A1(n6868), .A2(\mem[171][11] ), .B1(n6789), .B2(
        \mem[190][11] ), .ZN(n5179) );
  AOI22D0 U1382 ( .A1(n6977), .A2(\mem[161][11] ), .B1(n6995), .B2(
        \mem[151][11] ), .ZN(n5178) );
  ND4D0 U1383 ( .A1(n5181), .A2(n5180), .A3(n5179), .A4(n5178), .ZN(n5192) );
  AOI22D0 U1384 ( .A1(n6530), .A2(\mem[187][11] ), .B1(n6829), .B2(
        \mem[166][11] ), .ZN(n5185) );
  AOI22D0 U1385 ( .A1(n6954), .A2(\mem[138][11] ), .B1(n6828), .B2(
        \mem[184][11] ), .ZN(n5184) );
  AOI22D0 U1386 ( .A1(n6927), .A2(\mem[153][11] ), .B1(n6869), .B2(
        \mem[177][11] ), .ZN(n5183) );
  AOI22D0 U1387 ( .A1(n6525), .A2(\mem[163][11] ), .B1(n6733), .B2(
        \mem[186][11] ), .ZN(n5182) );
  ND4D0 U1388 ( .A1(n5185), .A2(n5184), .A3(n5183), .A4(n5182), .ZN(n5191) );
  AOI22D0 U1389 ( .A1(n6880), .A2(\mem[139][11] ), .B1(n6680), .B2(
        \mem[159][11] ), .ZN(n5189) );
  AOI22D0 U1390 ( .A1(n6819), .A2(\mem[189][11] ), .B1(n6901), .B2(
        \mem[137][11] ), .ZN(n5188) );
  AOI22D0 U1391 ( .A1(n6861), .A2(\mem[132][11] ), .B1(n6993), .B2(
        \mem[181][11] ), .ZN(n5187) );
  AOI22D0 U1392 ( .A1(n6979), .A2(\mem[142][11] ), .B1(n6882), .B2(
        \mem[143][11] ), .ZN(n5186) );
  ND4D0 U1393 ( .A1(n5189), .A2(n5188), .A3(n5187), .A4(n5186), .ZN(n5190) );
  NR4D0 U1394 ( .A1(n5193), .A2(n5192), .A3(n5191), .A4(n5190), .ZN(n5215) );
  AOI22D0 U1395 ( .A1(n6924), .A2(\mem[160][11] ), .B1(n6871), .B2(
        \mem[185][11] ), .ZN(n5197) );
  AOI22D0 U1396 ( .A1(n6953), .A2(\mem[175][11] ), .B1(n6174), .B2(
        \mem[182][11] ), .ZN(n5196) );
  AOI22D0 U1397 ( .A1(n6891), .A2(\mem[154][11] ), .B1(n6862), .B2(
        \mem[168][11] ), .ZN(n5195) );
  AOI22D0 U1398 ( .A1(n6981), .A2(\mem[188][11] ), .B1(n6698), .B2(
        \mem[130][11] ), .ZN(n5194) );
  ND4D0 U1399 ( .A1(n5197), .A2(n5196), .A3(n5195), .A4(n5194), .ZN(n5213) );
  AOI22D0 U1400 ( .A1(n6913), .A2(\mem[155][11] ), .B1(n6978), .B2(
        \mem[136][11] ), .ZN(n5200) );
  AOI22D0 U1401 ( .A1(n6784), .A2(\mem[156][11] ), .B1(n6922), .B2(
        \mem[157][11] ), .ZN(n5199) );
  AOI22D0 U1402 ( .A1(n6639), .A2(\mem[167][11] ), .B1(n6969), .B2(
        \mem[146][11] ), .ZN(n5198) );
  ND4D0 U1403 ( .A1(n5201), .A2(n5200), .A3(n5199), .A4(n5198), .ZN(n5212) );
  AOI22D0 U1404 ( .A1(n6658), .A2(\mem[178][11] ), .B1(n6988), .B2(
        \mem[191][11] ), .ZN(n5205) );
  AOI22D0 U1405 ( .A1(n6934), .A2(\mem[152][11] ), .B1(n6874), .B2(
        \mem[170][11] ), .ZN(n5204) );
  AOI22D0 U1406 ( .A1(n6890), .A2(\mem[164][11] ), .B1(n6906), .B2(
        \mem[140][11] ), .ZN(n5203) );
  AOI22D0 U1407 ( .A1(n6775), .A2(\mem[172][11] ), .B1(n6728), .B2(
        \mem[180][11] ), .ZN(n5202) );
  ND4D0 U1408 ( .A1(n5205), .A2(n5204), .A3(n5203), .A4(n5202), .ZN(n5211) );
  AOI22D0 U1409 ( .A1(n6830), .A2(\mem[135][11] ), .B1(n6923), .B2(
        \mem[162][11] ), .ZN(n5209) );
  AOI22D0 U1410 ( .A1(n6448), .A2(\mem[128][11] ), .B1(n6754), .B2(
        \mem[133][11] ), .ZN(n5208) );
  AOI22D0 U1411 ( .A1(n6916), .A2(\mem[149][11] ), .B1(n6964), .B2(
        \mem[158][11] ), .ZN(n5207) );
  AOI22D0 U1412 ( .A1(n6872), .A2(\mem[134][11] ), .B1(n6491), .B2(
        \mem[179][11] ), .ZN(n5206) );
  ND4D0 U1413 ( .A1(n5209), .A2(n5208), .A3(n5207), .A4(n5206), .ZN(n5210) );
  NR4D0 U1414 ( .A1(n5213), .A2(n5212), .A3(n5211), .A4(n5210), .ZN(n5214) );
  CKND2D0 U1415 ( .A1(n5215), .A2(n5214), .ZN(n5302) );
  AOI22D0 U1416 ( .A1(n6830), .A2(\mem[199][11] ), .B1(n6774), .B2(
        \mem[241][11] ), .ZN(n5219) );
  AOI22D0 U1417 ( .A1(n6727), .A2(\mem[234][11] ), .B1(n6923), .B2(
        \mem[226][11] ), .ZN(n5218) );
  AOI22D0 U1418 ( .A1(n6325), .A2(\mem[203][11] ), .B1(n6926), .B2(
        \mem[193][11] ), .ZN(n5217) );
  ND4D0 U1419 ( .A1(n5219), .A2(n5218), .A3(n5217), .A4(n5216), .ZN(n5235) );
  AOI22D0 U1420 ( .A1(n6881), .A2(\mem[208][11] ), .B1(n6902), .B2(
        \mem[229][11] ), .ZN(n5223) );
  AOI22D0 U1421 ( .A1(n6773), .A2(\mem[228][11] ), .B1(n6933), .B2(
        \mem[225][11] ), .ZN(n5222) );
  AOI22D0 U1422 ( .A1(n6917), .A2(\mem[238][11] ), .B1(n6639), .B2(
        \mem[231][11] ), .ZN(n5221) );
  AOI22D0 U1423 ( .A1(n6891), .A2(\mem[218][11] ), .B1(n6915), .B2(
        \mem[205][11] ), .ZN(n5220) );
  ND4D0 U1424 ( .A1(n5223), .A2(n5222), .A3(n5221), .A4(n5220), .ZN(n5234) );
  AOI22D0 U1425 ( .A1(n6747), .A2(\mem[212][11] ), .B1(n6889), .B2(
        \mem[220][11] ), .ZN(n5227) );
  AOI22D0 U1426 ( .A1(n6922), .A2(\mem[221][11] ), .B1(n6992), .B2(
        \mem[246][11] ), .ZN(n5226) );
  AOI22D0 U1427 ( .A1(n6791), .A2(\mem[224][11] ), .B1(n6982), .B2(
        \mem[194][11] ), .ZN(n5225) );
  AOI22D0 U1428 ( .A1(n6448), .A2(\mem[192][11] ), .B1(n6809), .B2(
        \mem[201][11] ), .ZN(n5224) );
  ND4D0 U1429 ( .A1(n5227), .A2(n5226), .A3(n5225), .A4(n5224), .ZN(n5233) );
  AOI22D0 U1430 ( .A1(n6802), .A2(\mem[216][11] ), .B1(n6979), .B2(
        \mem[206][11] ), .ZN(n5231) );
  AOI22D0 U1431 ( .A1(n6775), .A2(\mem[236][11] ), .B1(n6913), .B2(
        \mem[219][11] ), .ZN(n5230) );
  AOI22D0 U1432 ( .A1(n6907), .A2(\mem[195][11] ), .B1(n6863), .B2(
        \mem[247][11] ), .ZN(n5229) );
  AOI22D0 U1433 ( .A1(n6981), .A2(\mem[252][11] ), .B1(n6983), .B2(
        \mem[240][11] ), .ZN(n5228) );
  ND4D0 U1434 ( .A1(n5231), .A2(n5230), .A3(n5229), .A4(n5228), .ZN(n5232) );
  NR4D0 U1435 ( .A1(n5235), .A2(n5234), .A3(n5233), .A4(n5232), .ZN(n5257) );
  AOI22D0 U1436 ( .A1(n6835), .A2(\mem[196][11] ), .B1(n6837), .B2(
        \mem[207][11] ), .ZN(n5239) );
  AOI22D0 U1437 ( .A1(n6904), .A2(\mem[211][11] ), .B1(n6957), .B2(
        \mem[249][11] ), .ZN(n5238) );
  AOI22D0 U1438 ( .A1(n6955), .A2(\mem[213][11] ), .B1(n6912), .B2(
        \mem[248][11] ), .ZN(n5236) );
  ND4D0 U1439 ( .A1(n5239), .A2(n5238), .A3(n5237), .A4(n5236), .ZN(n5255) );
  AOI22D0 U1440 ( .A1(n6491), .A2(\mem[243][11] ), .B1(n6993), .B2(
        \mem[245][11] ), .ZN(n5243) );
  AOI22D0 U1441 ( .A1(n6995), .A2(\mem[215][11] ), .B1(n6990), .B2(
        \mem[204][11] ), .ZN(n5242) );
  AOI22D0 U1442 ( .A1(n6989), .A2(\mem[198][11] ), .B1(n6760), .B2(
        \mem[237][11] ), .ZN(n5241) );
  AOI22D0 U1443 ( .A1(n6868), .A2(\mem[235][11] ), .B1(n5966), .B2(
        \mem[223][11] ), .ZN(n5240) );
  ND4D0 U1444 ( .A1(n5243), .A2(n5242), .A3(n5241), .A4(n5240), .ZN(n5254) );
  AOI22D0 U1445 ( .A1(n6958), .A2(\mem[209][11] ), .B1(n6968), .B2(
        \mem[233][11] ), .ZN(n5247) );
  AOI22D0 U1446 ( .A1(n6733), .A2(\mem[250][11] ), .B1(n6994), .B2(
        \mem[254][11] ), .ZN(n5246) );
  AOI22D0 U1447 ( .A1(n6530), .A2(\mem[251][11] ), .B1(n6829), .B2(
        \mem[230][11] ), .ZN(n5245) );
  AOI22D0 U1448 ( .A1(n6525), .A2(\mem[227][11] ), .B1(n6873), .B2(
        \mem[222][11] ), .ZN(n5244) );
  AOI22D0 U1449 ( .A1(n6542), .A2(\mem[210][11] ), .B1(n6862), .B2(
        \mem[232][11] ), .ZN(n5251) );
  AOI22D0 U1450 ( .A1(n6819), .A2(\mem[253][11] ), .B1(n6935), .B2(
        \mem[255][11] ), .ZN(n5250) );
  AOI22D0 U1451 ( .A1(n6952), .A2(\mem[214][11] ), .B1(n6658), .B2(
        \mem[242][11] ), .ZN(n5249) );
  AOI22D0 U1452 ( .A1(n6179), .A2(\mem[239][11] ), .B1(n6954), .B2(
        \mem[202][11] ), .ZN(n5248) );
  ND4D0 U1453 ( .A1(n5251), .A2(n5250), .A3(n5249), .A4(n5248), .ZN(n5252) );
  NR4D0 U1454 ( .A1(n5255), .A2(n5254), .A3(n5253), .A4(n5252), .ZN(n5256) );
  AOI21D0 U1455 ( .A1(n5257), .A2(n5256), .B(n6945), .ZN(n5301) );
  AOI22D0 U1456 ( .A1(n6830), .A2(\mem[71][11] ), .B1(n6869), .B2(
        \mem[113][11] ), .ZN(n5261) );
  AOI22D0 U1457 ( .A1(n6829), .A2(\mem[102][11] ), .B1(n6863), .B2(
        \mem[119][11] ), .ZN(n5259) );
  AOI22D0 U1458 ( .A1(n6994), .A2(\mem[126][11] ), .B1(n6957), .B2(
        \mem[121][11] ), .ZN(n5258) );
  ND4D0 U1459 ( .A1(n5261), .A2(n5260), .A3(n5259), .A4(n5258), .ZN(n5277) );
  AOI22D0 U1460 ( .A1(n6861), .A2(\mem[68][11] ), .B1(n6658), .B2(
        \mem[114][11] ), .ZN(n5265) );
  AOI22D0 U1461 ( .A1(n6639), .A2(\mem[103][11] ), .B1(n6698), .B2(
        \mem[66][11] ), .ZN(n5264) );
  AOI22D0 U1462 ( .A1(n6775), .A2(\mem[108][11] ), .B1(n6842), .B2(
        \mem[90][11] ), .ZN(n5263) );
  AOI22D0 U1463 ( .A1(n6958), .A2(\mem[81][11] ), .B1(n6804), .B2(
        \mem[83][11] ), .ZN(n5262) );
  ND4D0 U1464 ( .A1(n5265), .A2(n5264), .A3(n5263), .A4(n5262), .ZN(n5276) );
  AOI22D0 U1465 ( .A1(n6868), .A2(\mem[107][11] ), .B1(n6923), .B2(
        \mem[98][11] ), .ZN(n5269) );
  AOI22D0 U1466 ( .A1(n6914), .A2(\mem[69][11] ), .B1(n6882), .B2(
        \mem[79][11] ), .ZN(n5268) );
  AOI22D0 U1467 ( .A1(n6880), .A2(\mem[75][11] ), .B1(n6955), .B2(
        \mem[85][11] ), .ZN(n5267) );
  AOI22D0 U1468 ( .A1(n6952), .A2(\mem[86][11] ), .B1(n6925), .B2(
        \mem[109][11] ), .ZN(n5266) );
  ND4D0 U1469 ( .A1(n5269), .A2(n5268), .A3(n5267), .A4(n5266), .ZN(n5275) );
  AOI22D0 U1470 ( .A1(n6847), .A2(\mem[89][11] ), .B1(n6988), .B2(
        \mem[127][11] ), .ZN(n5273) );
  AOI22D0 U1471 ( .A1(n6491), .A2(\mem[115][11] ), .B1(n6738), .B2(
        \mem[101][11] ), .ZN(n5272) );
  AOI22D0 U1472 ( .A1(n6448), .A2(\mem[64][11] ), .B1(n6992), .B2(
        \mem[118][11] ), .ZN(n5271) );
  AOI22D0 U1473 ( .A1(n6981), .A2(\mem[124][11] ), .B1(n6993), .B2(
        \mem[117][11] ), .ZN(n5270) );
  ND4D0 U1474 ( .A1(n5273), .A2(n5272), .A3(n5271), .A4(n5270), .ZN(n5274) );
  NR4D0 U1475 ( .A1(n5277), .A2(n5276), .A3(n5275), .A4(n5274), .ZN(n5299) );
  AOI22D0 U1476 ( .A1(n6728), .A2(\mem[116][11] ), .B1(n6968), .B2(
        \mem[105][11] ), .ZN(n5280) );
  AOI22D0 U1477 ( .A1(n6953), .A2(\mem[111][11] ), .B1(n6791), .B2(
        \mem[96][11] ), .ZN(n5279) );
  AOI22D0 U1478 ( .A1(n6934), .A2(\mem[88][11] ), .B1(n6959), .B2(
        \mem[67][11] ), .ZN(n5278) );
  ND4D0 U1479 ( .A1(n5281), .A2(n5280), .A3(n5279), .A4(n5278), .ZN(n5297) );
  AOI22D0 U1480 ( .A1(n6917), .A2(\mem[110][11] ), .B1(n6862), .B2(
        \mem[104][11] ), .ZN(n5285) );
  AOI22D0 U1481 ( .A1(n6954), .A2(\mem[74][11] ), .B1(n6828), .B2(
        \mem[120][11] ), .ZN(n5284) );
  AOI22D0 U1482 ( .A1(n6790), .A2(\mem[91][11] ), .B1(n6906), .B2(
        \mem[76][11] ), .ZN(n5283) );
  AOI22D0 U1483 ( .A1(n6819), .A2(\mem[125][11] ), .B1(n6542), .B2(
        \mem[82][11] ), .ZN(n5282) );
  ND4D0 U1484 ( .A1(n5285), .A2(n5284), .A3(n5283), .A4(n5282), .ZN(n5296) );
  AOI22D0 U1485 ( .A1(n6680), .A2(\mem[95][11] ), .B1(n6922), .B2(
        \mem[93][11] ), .ZN(n5289) );
  AOI22D0 U1486 ( .A1(n6881), .A2(\mem[80][11] ), .B1(n6733), .B2(
        \mem[122][11] ), .ZN(n5288) );
  AOI22D0 U1487 ( .A1(n6784), .A2(\mem[92][11] ), .B1(n6809), .B2(
        \mem[73][11] ), .ZN(n5287) );
  AOI22D0 U1488 ( .A1(n6727), .A2(\mem[106][11] ), .B1(n6964), .B2(
        \mem[94][11] ), .ZN(n5286) );
  ND4D0 U1489 ( .A1(n5289), .A2(n5288), .A3(n5287), .A4(n5286), .ZN(n5295) );
  AOI22D0 U1490 ( .A1(n6773), .A2(\mem[100][11] ), .B1(n6905), .B2(
        \mem[123][11] ), .ZN(n5293) );
  AOI22D0 U1491 ( .A1(n6747), .A2(\mem[84][11] ), .B1(n6978), .B2(
        \mem[72][11] ), .ZN(n5292) );
  AOI22D0 U1492 ( .A1(n6977), .A2(\mem[97][11] ), .B1(n6965), .B2(
        \mem[77][11] ), .ZN(n5291) );
  ND4D0 U1493 ( .A1(n5293), .A2(n5292), .A3(n5291), .A4(n5290), .ZN(n5294) );
  NR4D0 U1494 ( .A1(n5297), .A2(n5296), .A3(n5295), .A4(n5294), .ZN(n5298) );
  AOI21D0 U1495 ( .A1(n5299), .A2(n5298), .B(n7004), .ZN(n5300) );
  AOI211D0 U1496 ( .A1(n6951), .A2(n5302), .B(n5301), .C(n5300), .ZN(n5324) );
  AOI22D0 U1497 ( .A1(n6861), .A2(\mem[4][11] ), .B1(n6990), .B2(\mem[12][11] ), .ZN(n5306) );
  AOI22D0 U1498 ( .A1(n6773), .A2(\mem[36][11] ), .B1(n6892), .B2(
        \mem[44][11] ), .ZN(n5305) );
  AOI22D0 U1499 ( .A1(n6870), .A2(\mem[60][11] ), .B1(n6903), .B2(
        \mem[51][11] ), .ZN(n5304) );
  AOI22D0 U1500 ( .A1(n6993), .A2(\mem[53][11] ), .B1(n6916), .B2(
        \mem[21][11] ), .ZN(n5303) );
  ND4D0 U1501 ( .A1(n5306), .A2(n5305), .A3(n5304), .A4(n5303), .ZN(n5322) );
  AOI22D0 U1502 ( .A1(n6868), .A2(\mem[43][11] ), .B1(n6904), .B2(
        \mem[19][11] ), .ZN(n5310) );
  AOI22D0 U1503 ( .A1(n6830), .A2(\mem[7][11] ), .B1(n5966), .B2(\mem[31][11] ), .ZN(n5309) );
  AOI22D0 U1504 ( .A1(n6953), .A2(\mem[47][11] ), .B1(n6862), .B2(
        \mem[40][11] ), .ZN(n5307) );
  ND4D0 U1505 ( .A1(n5310), .A2(n5309), .A3(n5308), .A4(n5307), .ZN(n5321) );
  AOI22D0 U1506 ( .A1(n6952), .A2(\mem[22][11] ), .B1(n6880), .B2(
        \mem[11][11] ), .ZN(n5314) );
  AOI22D0 U1507 ( .A1(n6707), .A2(\mem[23][11] ), .B1(n6760), .B2(
        \mem[45][11] ), .ZN(n5313) );
  AOI22D0 U1508 ( .A1(n6530), .A2(\mem[59][11] ), .B1(n6658), .B2(
        \mem[50][11] ), .ZN(n5312) );
  AOI22D0 U1509 ( .A1(n6814), .A2(\mem[1][11] ), .B1(n6874), .B2(\mem[42][11] ), .ZN(n5311) );
  AOI22D0 U1510 ( .A1(n6971), .A2(\mem[38][11] ), .B1(n6954), .B2(
        \mem[10][11] ), .ZN(n5318) );
  AOI22D0 U1511 ( .A1(n6847), .A2(\mem[25][11] ), .B1(n6968), .B2(
        \mem[41][11] ), .ZN(n5317) );
  AOI22D0 U1512 ( .A1(n6958), .A2(\mem[17][11] ), .B1(n6698), .B2(\mem[2][11] ), .ZN(n5316) );
  AOI22D0 U1513 ( .A1(n6969), .A2(\mem[18][11] ), .B1(n6733), .B2(
        \mem[58][11] ), .ZN(n5315) );
  ND4D0 U1514 ( .A1(n5318), .A2(n5317), .A3(n5316), .A4(n5315), .ZN(n5319) );
  NR4D0 U1515 ( .A1(n5322), .A2(n5321), .A3(n5320), .A4(n5319), .ZN(n5323) );
  AOI32D0 U1516 ( .A1(n5325), .A2(n5324), .A3(n5323), .B1(n6856), .B2(n5324), 
        .ZN(dout[11]) );
  AOI22D0 U1517 ( .A1(n6892), .A2(\mem[44][5] ), .B1(n6971), .B2(\mem[38][5] ), 
        .ZN(n5329) );
  AOI22D0 U1518 ( .A1(n6914), .A2(\mem[5][5] ), .B1(n6491), .B2(\mem[51][5] ), 
        .ZN(n5327) );
  AOI22D0 U1519 ( .A1(n6870), .A2(\mem[60][5] ), .B1(n6835), .B2(\mem[4][5] ), 
        .ZN(n5326) );
  ND4D0 U1520 ( .A1(n5329), .A2(n5328), .A3(n5327), .A4(n5326), .ZN(n5345) );
  AOI22D0 U1521 ( .A1(n6979), .A2(\mem[14][5] ), .B1(n6296), .B2(\mem[29][5] ), 
        .ZN(n5333) );
  AOI22D0 U1522 ( .A1(n6916), .A2(\mem[21][5] ), .B1(n6869), .B2(\mem[49][5] ), 
        .ZN(n5332) );
  AOI22D0 U1523 ( .A1(n6968), .A2(\mem[41][5] ), .B1(n6862), .B2(\mem[40][5] ), 
        .ZN(n5331) );
  AOI22D0 U1524 ( .A1(n6784), .A2(\mem[28][5] ), .B1(n6913), .B2(\mem[27][5] ), 
        .ZN(n5330) );
  ND4D0 U1525 ( .A1(n5333), .A2(n5332), .A3(n5331), .A4(n5330), .ZN(n5344) );
  AOI22D0 U1526 ( .A1(n6977), .A2(\mem[33][5] ), .B1(n6658), .B2(\mem[50][5] ), 
        .ZN(n5337) );
  AOI22D0 U1527 ( .A1(n6912), .A2(\mem[56][5] ), .B1(n6990), .B2(\mem[12][5] ), 
        .ZN(n5336) );
  AOI22D0 U1528 ( .A1(n6749), .A2(\mem[43][5] ), .B1(n6957), .B2(\mem[57][5] ), 
        .ZN(n5335) );
  AOI22D0 U1529 ( .A1(n6928), .A2(\mem[7][5] ), .B1(n6863), .B2(\mem[55][5] ), 
        .ZN(n5334) );
  ND4D0 U1530 ( .A1(n5337), .A2(n5336), .A3(n5335), .A4(n5334), .ZN(n5343) );
  AOI22D0 U1531 ( .A1(n5966), .A2(\mem[31][5] ), .B1(n6707), .B2(\mem[23][5] ), 
        .ZN(n5341) );
  AOI22D0 U1532 ( .A1(n6179), .A2(\mem[47][5] ), .B1(n6923), .B2(\mem[34][5] ), 
        .ZN(n5340) );
  AOI22D0 U1533 ( .A1(n6325), .A2(\mem[11][5] ), .B1(n6760), .B2(\mem[45][5] ), 
        .ZN(n5339) );
  ND4D0 U1534 ( .A1(n5341), .A2(n5340), .A3(n5339), .A4(n5338), .ZN(n5342) );
  NR4D0 U1535 ( .A1(n5345), .A2(n5344), .A3(n5343), .A4(n5342), .ZN(n5497) );
  AOI22D0 U1536 ( .A1(n6889), .A2(\mem[156][5] ), .B1(n6955), .B2(
        \mem[149][5] ), .ZN(n5349) );
  AOI22D0 U1537 ( .A1(n6530), .A2(\mem[187][5] ), .B1(n6913), .B2(
        \mem[155][5] ), .ZN(n5348) );
  AOI22D0 U1538 ( .A1(n6980), .A2(\mem[189][5] ), .B1(n6967), .B2(
        \mem[167][5] ), .ZN(n5347) );
  AOI22D0 U1539 ( .A1(n6658), .A2(\mem[178][5] ), .B1(n6871), .B2(
        \mem[185][5] ), .ZN(n5346) );
  AOI22D0 U1540 ( .A1(n6934), .A2(\mem[152][5] ), .B1(n6979), .B2(
        \mem[142][5] ), .ZN(n5353) );
  AOI22D0 U1541 ( .A1(n6861), .A2(\mem[132][5] ), .B1(n6993), .B2(
        \mem[181][5] ), .ZN(n5351) );
  AOI22D0 U1542 ( .A1(n6879), .A2(\mem[186][5] ), .B1(n6837), .B2(
        \mem[143][5] ), .ZN(n5350) );
  ND4D0 U1543 ( .A1(n5353), .A2(n5352), .A3(n5351), .A4(n5350), .ZN(n5364) );
  AOI22D0 U1544 ( .A1(n6775), .A2(\mem[172][5] ), .B1(n6847), .B2(
        \mem[153][5] ), .ZN(n5357) );
  AOI22D0 U1545 ( .A1(n6958), .A2(\mem[145][5] ), .B1(n6906), .B2(
        \mem[140][5] ), .ZN(n5356) );
  AOI22D0 U1546 ( .A1(n6933), .A2(\mem[161][5] ), .B1(n6888), .B2(
        \mem[128][5] ), .ZN(n5355) );
  AOI22D0 U1547 ( .A1(n6969), .A2(\mem[146][5] ), .B1(n6296), .B2(
        \mem[157][5] ), .ZN(n5354) );
  ND4D0 U1548 ( .A1(n5357), .A2(n5356), .A3(n5355), .A4(n5354), .ZN(n5363) );
  AOI22D0 U1549 ( .A1(n6179), .A2(\mem[175][5] ), .B1(n6925), .B2(
        \mem[173][5] ), .ZN(n5361) );
  AOI22D0 U1550 ( .A1(n6325), .A2(\mem[139][5] ), .B1(n6814), .B2(
        \mem[129][5] ), .ZN(n5360) );
  AOI22D0 U1551 ( .A1(n6860), .A2(\mem[163][5] ), .B1(n6836), .B2(
        \mem[138][5] ), .ZN(n5359) );
  AOI22D0 U1552 ( .A1(n6859), .A2(\mem[180][5] ), .B1(n6964), .B2(
        \mem[158][5] ), .ZN(n5358) );
  ND4D0 U1553 ( .A1(n5361), .A2(n5360), .A3(n5359), .A4(n5358), .ZN(n5362) );
  NR4D0 U1554 ( .A1(n5365), .A2(n5364), .A3(n5363), .A4(n5362), .ZN(n5387) );
  AOI22D0 U1555 ( .A1(n6727), .A2(\mem[170][5] ), .B1(n6774), .B2(
        \mem[177][5] ), .ZN(n5369) );
  AOI22D0 U1556 ( .A1(n6935), .A2(\mem[191][5] ), .B1(n6956), .B2(
        \mem[168][5] ), .ZN(n5368) );
  AOI22D0 U1557 ( .A1(n6981), .A2(\mem[188][5] ), .B1(n6959), .B2(
        \mem[131][5] ), .ZN(n5367) );
  AOI22D0 U1558 ( .A1(n6614), .A2(\mem[150][5] ), .B1(n6991), .B2(
        \mem[148][5] ), .ZN(n5366) );
  ND4D0 U1559 ( .A1(n5369), .A2(n5368), .A3(n5367), .A4(n5366), .ZN(n5385) );
  AOI22D0 U1560 ( .A1(n6928), .A2(\mem[135][5] ), .B1(n6680), .B2(
        \mem[159][5] ), .ZN(n5372) );
  AOI22D0 U1561 ( .A1(n6995), .A2(\mem[151][5] ), .B1(n6968), .B2(
        \mem[169][5] ), .ZN(n5371) );
  AOI22D0 U1562 ( .A1(n6989), .A2(\mem[134][5] ), .B1(n6923), .B2(
        \mem[162][5] ), .ZN(n5370) );
  ND4D0 U1563 ( .A1(n5373), .A2(n5372), .A3(n5371), .A4(n5370), .ZN(n5384) );
  AOI22D0 U1564 ( .A1(n6983), .A2(\mem[176][5] ), .B1(n6891), .B2(
        \mem[154][5] ), .ZN(n5377) );
  AOI22D0 U1565 ( .A1(n6971), .A2(\mem[166][5] ), .B1(n6924), .B2(
        \mem[160][5] ), .ZN(n5376) );
  AOI22D0 U1566 ( .A1(n6901), .A2(\mem[137][5] ), .B1(n6903), .B2(
        \mem[179][5] ), .ZN(n5375) );
  AOI22D0 U1567 ( .A1(n6881), .A2(\mem[144][5] ), .B1(n6863), .B2(
        \mem[183][5] ), .ZN(n5374) );
  ND4D0 U1568 ( .A1(n5377), .A2(n5376), .A3(n5375), .A4(n5374), .ZN(n5383) );
  AOI22D0 U1569 ( .A1(n6982), .A2(\mem[130][5] ), .B1(n6828), .B2(
        \mem[184][5] ), .ZN(n5381) );
  AOI22D0 U1570 ( .A1(n6773), .A2(\mem[164][5] ), .B1(n6738), .B2(
        \mem[165][5] ), .ZN(n5380) );
  AOI22D0 U1571 ( .A1(n6994), .A2(\mem[190][5] ), .B1(n6174), .B2(
        \mem[182][5] ), .ZN(n5379) );
  AOI22D0 U1572 ( .A1(n6165), .A2(\mem[174][5] ), .B1(n6868), .B2(
        \mem[171][5] ), .ZN(n5378) );
  ND4D0 U1573 ( .A1(n5381), .A2(n5380), .A3(n5379), .A4(n5378), .ZN(n5382) );
  NR4D0 U1574 ( .A1(n5385), .A2(n5384), .A3(n5383), .A4(n5382), .ZN(n5386) );
  CKND2D0 U1575 ( .A1(n5387), .A2(n5386), .ZN(n5474) );
  AOI22D0 U1576 ( .A1(n6883), .A2(\mem[112][5] ), .B1(n6862), .B2(
        \mem[104][5] ), .ZN(n5391) );
  AOI22D0 U1577 ( .A1(n6525), .A2(\mem[99][5] ), .B1(n6728), .B2(\mem[116][5] ), .ZN(n5390) );
  AOI22D0 U1578 ( .A1(n6680), .A2(\mem[95][5] ), .B1(n6659), .B2(\mem[117][5] ), .ZN(n5389) );
  ND4D0 U1579 ( .A1(n5391), .A2(n5390), .A3(n5389), .A4(n5388), .ZN(n5407) );
  AOI22D0 U1580 ( .A1(n6836), .A2(\mem[74][5] ), .B1(n6968), .B2(\mem[105][5] ), .ZN(n5395) );
  AOI22D0 U1581 ( .A1(n6959), .A2(\mem[67][5] ), .B1(n6861), .B2(\mem[68][5] ), 
        .ZN(n5394) );
  AOI22D0 U1582 ( .A1(n6802), .A2(\mem[88][5] ), .B1(n6874), .B2(\mem[106][5] ), .ZN(n5393) );
  AOI22D0 U1583 ( .A1(n6325), .A2(\mem[75][5] ), .B1(n6863), .B2(\mem[119][5] ), .ZN(n5392) );
  ND4D0 U1584 ( .A1(n5395), .A2(n5394), .A3(n5393), .A4(n5392), .ZN(n5406) );
  AOI22D0 U1585 ( .A1(n6905), .A2(\mem[123][5] ), .B1(n6935), .B2(
        \mem[127][5] ), .ZN(n5399) );
  AOI22D0 U1586 ( .A1(n6707), .A2(\mem[87][5] ), .B1(n6869), .B2(\mem[113][5] ), .ZN(n5398) );
  AOI22D0 U1587 ( .A1(n6927), .A2(\mem[89][5] ), .B1(n6925), .B2(\mem[109][5] ), .ZN(n5397) );
  AOI22D0 U1588 ( .A1(n6892), .A2(\mem[108][5] ), .B1(n6842), .B2(\mem[90][5] ), .ZN(n5396) );
  ND4D0 U1589 ( .A1(n5399), .A2(n5398), .A3(n5397), .A4(n5396), .ZN(n5405) );
  AOI22D0 U1590 ( .A1(n6773), .A2(\mem[100][5] ), .B1(n6906), .B2(\mem[76][5] ), .ZN(n5403) );
  AOI22D0 U1591 ( .A1(n6913), .A2(\mem[91][5] ), .B1(n6698), .B2(\mem[66][5] ), 
        .ZN(n5402) );
  AOI22D0 U1592 ( .A1(n6903), .A2(\mem[115][5] ), .B1(n6174), .B2(
        \mem[118][5] ), .ZN(n5401) );
  AOI22D0 U1593 ( .A1(n6957), .A2(\mem[121][5] ), .B1(n6837), .B2(\mem[79][5] ), .ZN(n5400) );
  ND4D0 U1594 ( .A1(n5403), .A2(n5402), .A3(n5401), .A4(n5400), .ZN(n5404) );
  NR4D0 U1595 ( .A1(n5407), .A2(n5406), .A3(n5405), .A4(n5404), .ZN(n5429) );
  AOI22D0 U1596 ( .A1(n6784), .A2(\mem[92][5] ), .B1(n6923), .B2(\mem[98][5] ), 
        .ZN(n5411) );
  AOI22D0 U1597 ( .A1(n6749), .A2(\mem[107][5] ), .B1(n6915), .B2(\mem[77][5] ), .ZN(n5410) );
  AOI22D0 U1598 ( .A1(n6614), .A2(\mem[86][5] ), .B1(n6916), .B2(\mem[85][5] ), 
        .ZN(n5408) );
  ND4D0 U1599 ( .A1(n5411), .A2(n5410), .A3(n5409), .A4(n5408), .ZN(n5427) );
  AOI22D0 U1600 ( .A1(n6981), .A2(\mem[124][5] ), .B1(n6804), .B2(\mem[83][5] ), .ZN(n5415) );
  AOI22D0 U1601 ( .A1(n6979), .A2(\mem[78][5] ), .B1(n6936), .B2(\mem[81][5] ), 
        .ZN(n5414) );
  AOI22D0 U1602 ( .A1(n6754), .A2(\mem[69][5] ), .B1(n6901), .B2(\mem[73][5] ), 
        .ZN(n5413) );
  AOI22D0 U1603 ( .A1(n6830), .A2(\mem[71][5] ), .B1(n6912), .B2(\mem[120][5] ), .ZN(n5412) );
  ND4D0 U1604 ( .A1(n5415), .A2(n5414), .A3(n5413), .A4(n5412), .ZN(n5426) );
  AOI22D0 U1605 ( .A1(n6179), .A2(\mem[111][5] ), .B1(n6296), .B2(\mem[93][5] ), .ZN(n5419) );
  AOI22D0 U1606 ( .A1(n6969), .A2(\mem[82][5] ), .B1(n6978), .B2(\mem[72][5] ), 
        .ZN(n5418) );
  AOI22D0 U1607 ( .A1(n6980), .A2(\mem[125][5] ), .B1(n6902), .B2(
        \mem[101][5] ), .ZN(n5417) );
  AOI22D0 U1608 ( .A1(n6926), .A2(\mem[65][5] ), .B1(n6991), .B2(\mem[84][5] ), 
        .ZN(n5416) );
  ND4D0 U1609 ( .A1(n5419), .A2(n5418), .A3(n5417), .A4(n5416), .ZN(n5425) );
  AOI22D0 U1610 ( .A1(n6989), .A2(\mem[70][5] ), .B1(n6967), .B2(\mem[103][5] ), .ZN(n5423) );
  AOI22D0 U1611 ( .A1(n6933), .A2(\mem[97][5] ), .B1(n6658), .B2(\mem[114][5] ), .ZN(n5422) );
  AOI22D0 U1612 ( .A1(n6879), .A2(\mem[122][5] ), .B1(n6789), .B2(
        \mem[126][5] ), .ZN(n5421) );
  AOI22D0 U1613 ( .A1(n6970), .A2(\mem[80][5] ), .B1(n6888), .B2(\mem[64][5] ), 
        .ZN(n5420) );
  NR4D0 U1614 ( .A1(n5427), .A2(n5426), .A3(n5425), .A4(n5424), .ZN(n5428) );
  AOI22D0 U1615 ( .A1(n6819), .A2(\mem[253][5] ), .B1(n6991), .B2(
        \mem[212][5] ), .ZN(n5433) );
  AOI22D0 U1616 ( .A1(n6905), .A2(\mem[251][5] ), .B1(n6738), .B2(
        \mem[229][5] ), .ZN(n5431) );
  AOI22D0 U1617 ( .A1(n6863), .A2(\mem[247][5] ), .B1(n6994), .B2(
        \mem[254][5] ), .ZN(n5430) );
  ND4D0 U1618 ( .A1(n5433), .A2(n5432), .A3(n5431), .A4(n5430), .ZN(n5449) );
  AOI22D0 U1619 ( .A1(n6165), .A2(\mem[238][5] ), .B1(n6861), .B2(
        \mem[196][5] ), .ZN(n5437) );
  AOI22D0 U1620 ( .A1(n6890), .A2(\mem[228][5] ), .B1(n6969), .B2(
        \mem[210][5] ), .ZN(n5436) );
  AOI22D0 U1621 ( .A1(n6680), .A2(\mem[223][5] ), .B1(n6966), .B2(
        \mem[242][5] ), .ZN(n5435) );
  AOI22D0 U1622 ( .A1(n6993), .A2(\mem[245][5] ), .B1(n6174), .B2(
        \mem[246][5] ), .ZN(n5434) );
  ND4D0 U1623 ( .A1(n5437), .A2(n5436), .A3(n5435), .A4(n5434), .ZN(n5448) );
  AOI22D0 U1624 ( .A1(n6879), .A2(\mem[250][5] ), .B1(n6874), .B2(
        \mem[234][5] ), .ZN(n5441) );
  AOI22D0 U1625 ( .A1(n6790), .A2(\mem[219][5] ), .B1(n6828), .B2(
        \mem[248][5] ), .ZN(n5440) );
  AOI22D0 U1626 ( .A1(n6842), .A2(\mem[218][5] ), .B1(n6925), .B2(
        \mem[237][5] ), .ZN(n5439) );
  AOI22D0 U1627 ( .A1(n6958), .A2(\mem[209][5] ), .B1(n6563), .B2(
        \mem[200][5] ), .ZN(n5438) );
  ND4D0 U1628 ( .A1(n5441), .A2(n5440), .A3(n5439), .A4(n5438), .ZN(n5447) );
  AOI22D0 U1629 ( .A1(n6926), .A2(\mem[193][5] ), .B1(n6957), .B2(
        \mem[249][5] ), .ZN(n5445) );
  AOI22D0 U1630 ( .A1(n6614), .A2(\mem[214][5] ), .B1(n6754), .B2(
        \mem[197][5] ), .ZN(n5444) );
  AOI22D0 U1631 ( .A1(n6971), .A2(\mem[230][5] ), .B1(n6935), .B2(
        \mem[255][5] ), .ZN(n5443) );
  AOI22D0 U1632 ( .A1(n6870), .A2(\mem[252][5] ), .B1(n6707), .B2(
        \mem[215][5] ), .ZN(n5442) );
  ND4D0 U1633 ( .A1(n5445), .A2(n5444), .A3(n5443), .A4(n5442), .ZN(n5446) );
  NR4D0 U1634 ( .A1(n5449), .A2(n5448), .A3(n5447), .A4(n5446), .ZN(n5471) );
  AOI22D0 U1635 ( .A1(n6983), .A2(\mem[240][5] ), .B1(n6859), .B2(
        \mem[244][5] ), .ZN(n5452) );
  AOI22D0 U1636 ( .A1(n6955), .A2(\mem[213][5] ), .B1(n6837), .B2(
        \mem[207][5] ), .ZN(n5451) );
  AOI22D0 U1637 ( .A1(n6959), .A2(\mem[195][5] ), .B1(n6903), .B2(
        \mem[243][5] ), .ZN(n5450) );
  ND4D0 U1638 ( .A1(n5453), .A2(n5452), .A3(n5451), .A4(n5450), .ZN(n5469) );
  AOI22D0 U1639 ( .A1(n6639), .A2(\mem[231][5] ), .B1(n6923), .B2(
        \mem[226][5] ), .ZN(n5457) );
  AOI22D0 U1640 ( .A1(n6448), .A2(\mem[192][5] ), .B1(n6965), .B2(
        \mem[205][5] ), .ZN(n5456) );
  AOI22D0 U1641 ( .A1(n6296), .A2(\mem[221][5] ), .B1(n6804), .B2(
        \mem[211][5] ), .ZN(n5455) );
  AOI22D0 U1642 ( .A1(n6892), .A2(\mem[236][5] ), .B1(n6748), .B2(
        \mem[233][5] ), .ZN(n5454) );
  ND4D0 U1643 ( .A1(n5457), .A2(n5456), .A3(n5455), .A4(n5454), .ZN(n5468) );
  AOI22D0 U1644 ( .A1(n6954), .A2(\mem[202][5] ), .B1(n6982), .B2(
        \mem[194][5] ), .ZN(n5461) );
  AOI22D0 U1645 ( .A1(n6970), .A2(\mem[208][5] ), .B1(n6906), .B2(
        \mem[204][5] ), .ZN(n5460) );
  AOI22D0 U1646 ( .A1(n6749), .A2(\mem[235][5] ), .B1(n6989), .B2(
        \mem[198][5] ), .ZN(n5459) );
  AOI22D0 U1647 ( .A1(n6860), .A2(\mem[227][5] ), .B1(n6809), .B2(
        \mem[201][5] ), .ZN(n5458) );
  ND4D0 U1648 ( .A1(n5461), .A2(n5460), .A3(n5459), .A4(n5458), .ZN(n5467) );
  AOI22D0 U1649 ( .A1(n6933), .A2(\mem[225][5] ), .B1(n6924), .B2(
        \mem[224][5] ), .ZN(n5465) );
  AOI22D0 U1650 ( .A1(n6862), .A2(\mem[232][5] ), .B1(n6964), .B2(
        \mem[222][5] ), .ZN(n5464) );
  AOI22D0 U1651 ( .A1(n6759), .A2(\mem[206][5] ), .B1(n6889), .B2(
        \mem[220][5] ), .ZN(n5463) );
  ND4D0 U1652 ( .A1(n5465), .A2(n5464), .A3(n5463), .A4(n5462), .ZN(n5466) );
  NR4D0 U1653 ( .A1(n5469), .A2(n5468), .A3(n5467), .A4(n5466), .ZN(n5470) );
  AOI21D0 U1654 ( .A1(n5471), .A2(n5470), .B(n6945), .ZN(n5472) );
  AOI22D0 U1655 ( .A1(n6728), .A2(\mem[52][5] ), .B1(n6936), .B2(\mem[17][5] ), 
        .ZN(n5478) );
  AOI22D0 U1656 ( .A1(n6860), .A2(\mem[35][5] ), .B1(n6902), .B2(\mem[37][5] ), 
        .ZN(n5477) );
  AOI22D0 U1657 ( .A1(n6872), .A2(\mem[6][5] ), .B1(n6789), .B2(\mem[62][5] ), 
        .ZN(n5476) );
  AOI22D0 U1658 ( .A1(n6890), .A2(\mem[36][5] ), .B1(n6873), .B2(\mem[30][5] ), 
        .ZN(n5475) );
  ND4D0 U1659 ( .A1(n5478), .A2(n5477), .A3(n5476), .A4(n5475), .ZN(n5494) );
  AOI22D0 U1660 ( .A1(n6791), .A2(\mem[32][5] ), .B1(n6563), .B2(\mem[8][5] ), 
        .ZN(n5482) );
  AOI22D0 U1661 ( .A1(n6959), .A2(\mem[3][5] ), .B1(n6698), .B2(\mem[2][5] ), 
        .ZN(n5481) );
  AOI22D0 U1662 ( .A1(n6614), .A2(\mem[22][5] ), .B1(n6847), .B2(\mem[25][5] ), 
        .ZN(n5480) );
  AOI22D0 U1663 ( .A1(n6814), .A2(\mem[1][5] ), .B1(n6988), .B2(\mem[63][5] ), 
        .ZN(n5479) );
  ND4D0 U1664 ( .A1(n5482), .A2(n5481), .A3(n5480), .A4(n5479), .ZN(n5493) );
  AOI22D0 U1665 ( .A1(n6165), .A2(\mem[46][5] ), .B1(n6804), .B2(\mem[19][5] ), 
        .ZN(n5486) );
  AOI22D0 U1666 ( .A1(n6888), .A2(\mem[0][5] ), .B1(n6659), .B2(\mem[53][5] ), 
        .ZN(n5484) );
  AOI22D0 U1667 ( .A1(n6905), .A2(\mem[59][5] ), .B1(n6883), .B2(\mem[48][5] ), 
        .ZN(n5483) );
  ND4D0 U1668 ( .A1(n5486), .A2(n5485), .A3(n5484), .A4(n5483), .ZN(n5492) );
  AOI22D0 U1669 ( .A1(n6970), .A2(\mem[16][5] ), .B1(n6965), .B2(\mem[13][5] ), 
        .ZN(n5490) );
  AOI22D0 U1670 ( .A1(n6980), .A2(\mem[61][5] ), .B1(n6891), .B2(\mem[26][5] ), 
        .ZN(n5489) );
  AOI22D0 U1671 ( .A1(n6809), .A2(\mem[9][5] ), .B1(n6874), .B2(\mem[42][5] ), 
        .ZN(n5488) );
  AOI22D0 U1672 ( .A1(n6802), .A2(\mem[24][5] ), .B1(n6542), .B2(\mem[18][5] ), 
        .ZN(n5487) );
  ND4D0 U1673 ( .A1(n5490), .A2(n5489), .A3(n5488), .A4(n5487), .ZN(n5491) );
  NR4D0 U1674 ( .A1(n5494), .A2(n5493), .A3(n5492), .A4(n5491), .ZN(n5495) );
  AOI32D0 U1675 ( .A1(n5497), .A2(n5496), .A3(n5495), .B1(n6856), .B2(n5496), 
        .ZN(dout[5]) );
  AOI22D0 U1676 ( .A1(n6873), .A2(\mem[30][8] ), .B1(n6912), .B2(\mem[56][8] ), 
        .ZN(n5500) );
  AOI22D0 U1677 ( .A1(n6888), .A2(\mem[0][8] ), .B1(n6760), .B2(\mem[45][8] ), 
        .ZN(n5499) );
  AOI22D0 U1678 ( .A1(n6803), .A2(\mem[55][8] ), .B1(n6698), .B2(\mem[2][8] ), 
        .ZN(n5498) );
  ND4D0 U1679 ( .A1(n5501), .A2(n5500), .A3(n5499), .A4(n5498), .ZN(n5517) );
  AOI22D0 U1680 ( .A1(n6977), .A2(\mem[33][8] ), .B1(n6707), .B2(\mem[23][8] ), 
        .ZN(n5505) );
  AOI22D0 U1681 ( .A1(n6814), .A2(\mem[1][8] ), .B1(n6991), .B2(\mem[20][8] ), 
        .ZN(n5504) );
  AOI22D0 U1682 ( .A1(n6979), .A2(\mem[14][8] ), .B1(n6784), .B2(\mem[28][8] ), 
        .ZN(n5503) );
  AOI22D0 U1683 ( .A1(n6917), .A2(\mem[46][8] ), .B1(n6993), .B2(\mem[53][8] ), 
        .ZN(n5502) );
  ND4D0 U1684 ( .A1(n5505), .A2(n5504), .A3(n5503), .A4(n5502), .ZN(n5516) );
  AOI22D0 U1685 ( .A1(n6969), .A2(\mem[18][8] ), .B1(n6994), .B2(\mem[62][8] ), 
        .ZN(n5509) );
  AOI22D0 U1686 ( .A1(n6749), .A2(\mem[43][8] ), .B1(n6956), .B2(\mem[40][8] ), 
        .ZN(n5508) );
  AOI22D0 U1687 ( .A1(n6927), .A2(\mem[25][8] ), .B1(n6902), .B2(\mem[37][8] ), 
        .ZN(n5507) );
  AOI22D0 U1688 ( .A1(n6928), .A2(\mem[7][8] ), .B1(n6980), .B2(\mem[61][8] ), 
        .ZN(n5506) );
  ND4D0 U1689 ( .A1(n5509), .A2(n5508), .A3(n5507), .A4(n5506), .ZN(n5515) );
  AOI22D0 U1690 ( .A1(n6891), .A2(\mem[26][8] ), .B1(n6809), .B2(\mem[9][8] ), 
        .ZN(n5513) );
  AOI22D0 U1691 ( .A1(n6791), .A2(\mem[32][8] ), .B1(n6871), .B2(\mem[57][8] ), 
        .ZN(n5512) );
  AOI22D0 U1692 ( .A1(n6880), .A2(\mem[11][8] ), .B1(n6836), .B2(\mem[10][8] ), 
        .ZN(n5511) );
  ND4D0 U1693 ( .A1(n5513), .A2(n5512), .A3(n5511), .A4(n5510), .ZN(n5514) );
  NR4D0 U1694 ( .A1(n5517), .A2(n5516), .A3(n5515), .A4(n5514), .ZN(n5669) );
  AOI22D0 U1695 ( .A1(n6916), .A2(\mem[149][8] ), .B1(n6873), .B2(
        \mem[158][8] ), .ZN(n5521) );
  AOI22D0 U1696 ( .A1(n6905), .A2(\mem[187][8] ), .B1(n6989), .B2(
        \mem[134][8] ), .ZN(n5520) );
  AOI22D0 U1697 ( .A1(n6981), .A2(\mem[188][8] ), .B1(n6891), .B2(
        \mem[154][8] ), .ZN(n5519) );
  AOI22D0 U1698 ( .A1(n6835), .A2(\mem[132][8] ), .B1(n6728), .B2(
        \mem[180][8] ), .ZN(n5518) );
  ND4D0 U1699 ( .A1(n5521), .A2(n5520), .A3(n5519), .A4(n5518), .ZN(n5537) );
  AOI22D0 U1700 ( .A1(n6928), .A2(\mem[135][8] ), .B1(n6880), .B2(
        \mem[139][8] ), .ZN(n5525) );
  AOI22D0 U1701 ( .A1(n6902), .A2(\mem[165][8] ), .B1(n6882), .B2(
        \mem[143][8] ), .ZN(n5524) );
  AOI22D0 U1702 ( .A1(n6868), .A2(\mem[171][8] ), .B1(n6990), .B2(
        \mem[140][8] ), .ZN(n5523) );
  AOI22D0 U1703 ( .A1(n6959), .A2(\mem[131][8] ), .B1(n6862), .B2(
        \mem[168][8] ), .ZN(n5522) );
  ND4D0 U1704 ( .A1(n5525), .A2(n5524), .A3(n5523), .A4(n5522), .ZN(n5536) );
  AOI22D0 U1705 ( .A1(n6953), .A2(\mem[175][8] ), .B1(n6888), .B2(
        \mem[128][8] ), .ZN(n5529) );
  AOI22D0 U1706 ( .A1(n6991), .A2(\mem[148][8] ), .B1(n6863), .B2(
        \mem[183][8] ), .ZN(n5528) );
  AOI22D0 U1707 ( .A1(n6165), .A2(\mem[174][8] ), .B1(n6847), .B2(
        \mem[153][8] ), .ZN(n5527) );
  AOI22D0 U1708 ( .A1(n6933), .A2(\mem[161][8] ), .B1(n6965), .B2(
        \mem[141][8] ), .ZN(n5526) );
  ND4D0 U1709 ( .A1(n5529), .A2(n5528), .A3(n5527), .A4(n5526), .ZN(n5535) );
  AOI22D0 U1710 ( .A1(n6860), .A2(\mem[163][8] ), .B1(n6754), .B2(
        \mem[133][8] ), .ZN(n5533) );
  AOI22D0 U1711 ( .A1(n6922), .A2(\mem[157][8] ), .B1(n6912), .B2(
        \mem[184][8] ), .ZN(n5532) );
  AOI22D0 U1712 ( .A1(n6892), .A2(\mem[172][8] ), .B1(n6881), .B2(
        \mem[144][8] ), .ZN(n5530) );
  ND4D0 U1713 ( .A1(n5533), .A2(n5532), .A3(n5531), .A4(n5530), .ZN(n5534) );
  NR4D0 U1714 ( .A1(n5537), .A2(n5536), .A3(n5535), .A4(n5534), .ZN(n5559) );
  AOI22D0 U1715 ( .A1(n6924), .A2(\mem[160][8] ), .B1(n6982), .B2(
        \mem[130][8] ), .ZN(n5541) );
  AOI22D0 U1716 ( .A1(n6790), .A2(\mem[155][8] ), .B1(n6954), .B2(
        \mem[138][8] ), .ZN(n5540) );
  AOI22D0 U1717 ( .A1(n6952), .A2(\mem[150][8] ), .B1(n6925), .B2(
        \mem[173][8] ), .ZN(n5539) );
  AOI22D0 U1718 ( .A1(n6980), .A2(\mem[189][8] ), .B1(n6994), .B2(
        \mem[190][8] ), .ZN(n5538) );
  ND4D0 U1719 ( .A1(n5541), .A2(n5540), .A3(n5539), .A4(n5538), .ZN(n5557) );
  AOI22D0 U1720 ( .A1(n6890), .A2(\mem[164][8] ), .B1(n6968), .B2(
        \mem[169][8] ), .ZN(n5545) );
  AOI22D0 U1721 ( .A1(n6542), .A2(\mem[146][8] ), .B1(n6809), .B2(
        \mem[137][8] ), .ZN(n5544) );
  AOI22D0 U1722 ( .A1(n6879), .A2(\mem[186][8] ), .B1(n5966), .B2(
        \mem[159][8] ), .ZN(n5543) );
  AOI22D0 U1723 ( .A1(n6659), .A2(\mem[181][8] ), .B1(n6904), .B2(
        \mem[147][8] ), .ZN(n5542) );
  AOI22D0 U1724 ( .A1(n6814), .A2(\mem[129][8] ), .B1(n6966), .B2(
        \mem[178][8] ), .ZN(n5549) );
  AOI22D0 U1725 ( .A1(n6923), .A2(\mem[162][8] ), .B1(n6988), .B2(
        \mem[191][8] ), .ZN(n5548) );
  AOI22D0 U1726 ( .A1(n6869), .A2(\mem[177][8] ), .B1(n6992), .B2(
        \mem[182][8] ), .ZN(n5547) );
  AOI22D0 U1727 ( .A1(n6883), .A2(\mem[176][8] ), .B1(n6958), .B2(
        \mem[145][8] ), .ZN(n5546) );
  ND4D0 U1728 ( .A1(n5549), .A2(n5548), .A3(n5547), .A4(n5546), .ZN(n5555) );
  AOI22D0 U1729 ( .A1(n6971), .A2(\mem[166][8] ), .B1(n6903), .B2(
        \mem[179][8] ), .ZN(n5553) );
  AOI22D0 U1730 ( .A1(n6967), .A2(\mem[167][8] ), .B1(n6727), .B2(
        \mem[170][8] ), .ZN(n5551) );
  AOI22D0 U1731 ( .A1(n6802), .A2(\mem[152][8] ), .B1(n6979), .B2(
        \mem[142][8] ), .ZN(n5550) );
  ND4D0 U1732 ( .A1(n5553), .A2(n5552), .A3(n5551), .A4(n5550), .ZN(n5554) );
  NR4D0 U1733 ( .A1(n5557), .A2(n5556), .A3(n5555), .A4(n5554), .ZN(n5558) );
  CKND2D0 U1734 ( .A1(n5559), .A2(n5558), .ZN(n5646) );
  AOI22D0 U1735 ( .A1(n6179), .A2(\mem[239][8] ), .B1(n6835), .B2(
        \mem[196][8] ), .ZN(n5563) );
  AOI22D0 U1736 ( .A1(n6814), .A2(\mem[193][8] ), .B1(n6829), .B2(
        \mem[230][8] ), .ZN(n5562) );
  AOI22D0 U1737 ( .A1(n6979), .A2(\mem[206][8] ), .B1(n6880), .B2(
        \mem[203][8] ), .ZN(n5561) );
  AOI22D0 U1738 ( .A1(n6905), .A2(\mem[251][8] ), .B1(n6847), .B2(
        \mem[217][8] ), .ZN(n5560) );
  ND4D0 U1739 ( .A1(n5563), .A2(n5562), .A3(n5561), .A4(n5560), .ZN(n5579) );
  AOI22D0 U1740 ( .A1(n6868), .A2(\mem[235][8] ), .B1(n6924), .B2(
        \mem[224][8] ), .ZN(n5567) );
  AOI22D0 U1741 ( .A1(n6954), .A2(\mem[202][8] ), .B1(n6862), .B2(
        \mem[232][8] ), .ZN(n5566) );
  AOI22D0 U1742 ( .A1(n6959), .A2(\mem[195][8] ), .B1(n6707), .B2(
        \mem[215][8] ), .ZN(n5565) );
  AOI22D0 U1743 ( .A1(n6917), .A2(\mem[238][8] ), .B1(n6658), .B2(
        \mem[242][8] ), .ZN(n5564) );
  ND4D0 U1744 ( .A1(n5567), .A2(n5566), .A3(n5565), .A4(n5564), .ZN(n5578) );
  AOI22D0 U1745 ( .A1(n6863), .A2(\mem[247][8] ), .B1(n6728), .B2(
        \mem[244][8] ), .ZN(n5571) );
  AOI22D0 U1746 ( .A1(n6991), .A2(\mem[212][8] ), .B1(n6994), .B2(
        \mem[254][8] ), .ZN(n5570) );
  AOI22D0 U1747 ( .A1(n6860), .A2(\mem[227][8] ), .B1(n6925), .B2(
        \mem[237][8] ), .ZN(n5569) );
  AOI22D0 U1748 ( .A1(n6980), .A2(\mem[253][8] ), .B1(n6955), .B2(
        \mem[213][8] ), .ZN(n5568) );
  ND4D0 U1749 ( .A1(n5571), .A2(n5570), .A3(n5569), .A4(n5568), .ZN(n5577) );
  AOI22D0 U1750 ( .A1(n6659), .A2(\mem[245][8] ), .B1(n6958), .B2(
        \mem[209][8] ), .ZN(n5574) );
  AOI22D0 U1751 ( .A1(n6892), .A2(\mem[236][8] ), .B1(n6883), .B2(
        \mem[240][8] ), .ZN(n5573) );
  AOI22D0 U1752 ( .A1(n6968), .A2(\mem[233][8] ), .B1(n6912), .B2(
        \mem[248][8] ), .ZN(n5572) );
  ND4D0 U1753 ( .A1(n5575), .A2(n5574), .A3(n5573), .A4(n5572), .ZN(n5576) );
  NR4D0 U1754 ( .A1(n5579), .A2(n5578), .A3(n5577), .A4(n5576), .ZN(n5601) );
  AOI22D0 U1755 ( .A1(n6977), .A2(\mem[225][8] ), .B1(n6888), .B2(
        \mem[192][8] ), .ZN(n5583) );
  AOI22D0 U1756 ( .A1(n6989), .A2(\mem[198][8] ), .B1(n6491), .B2(
        \mem[243][8] ), .ZN(n5582) );
  AOI22D0 U1757 ( .A1(n6890), .A2(\mem[228][8] ), .B1(n6842), .B2(
        \mem[218][8] ), .ZN(n5581) );
  AOI22D0 U1758 ( .A1(n6969), .A2(\mem[210][8] ), .B1(n6923), .B2(
        \mem[226][8] ), .ZN(n5580) );
  ND4D0 U1759 ( .A1(n5583), .A2(n5582), .A3(n5581), .A4(n5580), .ZN(n5599) );
  AOI22D0 U1760 ( .A1(n6809), .A2(\mem[201][8] ), .B1(n6727), .B2(
        \mem[234][8] ), .ZN(n5587) );
  AOI22D0 U1761 ( .A1(n6680), .A2(\mem[223][8] ), .B1(n6837), .B2(
        \mem[207][8] ), .ZN(n5586) );
  AOI22D0 U1762 ( .A1(n6904), .A2(\mem[211][8] ), .B1(n6982), .B2(
        \mem[194][8] ), .ZN(n5585) );
  AOI22D0 U1763 ( .A1(n6296), .A2(\mem[221][8] ), .B1(n6871), .B2(
        \mem[249][8] ), .ZN(n5584) );
  ND4D0 U1764 ( .A1(n5587), .A2(n5586), .A3(n5585), .A4(n5584), .ZN(n5598) );
  AOI22D0 U1765 ( .A1(n6563), .A2(\mem[200][8] ), .B1(n6990), .B2(
        \mem[204][8] ), .ZN(n5591) );
  AOI22D0 U1766 ( .A1(n6935), .A2(\mem[255][8] ), .B1(n6873), .B2(
        \mem[222][8] ), .ZN(n5590) );
  AOI22D0 U1767 ( .A1(n6928), .A2(\mem[199][8] ), .B1(n6952), .B2(
        \mem[214][8] ), .ZN(n5589) );
  ND4D0 U1768 ( .A1(n5591), .A2(n5590), .A3(n5589), .A4(n5588), .ZN(n5597) );
  AOI22D0 U1769 ( .A1(n6870), .A2(\mem[252][8] ), .B1(n6733), .B2(
        \mem[250][8] ), .ZN(n5595) );
  AOI22D0 U1770 ( .A1(n6967), .A2(\mem[231][8] ), .B1(n6970), .B2(
        \mem[208][8] ), .ZN(n5594) );
  AOI22D0 U1771 ( .A1(n6889), .A2(\mem[220][8] ), .B1(n6869), .B2(
        \mem[241][8] ), .ZN(n5593) );
  AOI22D0 U1772 ( .A1(n6934), .A2(\mem[216][8] ), .B1(n6754), .B2(
        \mem[197][8] ), .ZN(n5592) );
  ND4D0 U1773 ( .A1(n5595), .A2(n5594), .A3(n5593), .A4(n5592), .ZN(n5596) );
  NR4D0 U1774 ( .A1(n5599), .A2(n5598), .A3(n5597), .A4(n5596), .ZN(n5600) );
  AOI21D0 U1775 ( .A1(n5601), .A2(n5600), .B(n6945), .ZN(n5645) );
  AOI22D0 U1776 ( .A1(n6913), .A2(\mem[91][8] ), .B1(n6904), .B2(\mem[83][8] ), 
        .ZN(n5605) );
  AOI22D0 U1777 ( .A1(n6881), .A2(\mem[80][8] ), .B1(n5966), .B2(\mem[95][8] ), 
        .ZN(n5604) );
  AOI22D0 U1778 ( .A1(n6979), .A2(\mem[78][8] ), .B1(n6955), .B2(\mem[85][8] ), 
        .ZN(n5603) );
  AOI22D0 U1779 ( .A1(n6953), .A2(\mem[111][8] ), .B1(n6614), .B2(\mem[86][8] ), .ZN(n5602) );
  ND4D0 U1780 ( .A1(n5605), .A2(n5604), .A3(n5603), .A4(n5602), .ZN(n5621) );
  AOI22D0 U1781 ( .A1(n6880), .A2(\mem[75][8] ), .B1(n6863), .B2(\mem[119][8] ), .ZN(n5609) );
  AOI22D0 U1782 ( .A1(n6922), .A2(\mem[93][8] ), .B1(n6995), .B2(\mem[87][8] ), 
        .ZN(n5608) );
  AOI22D0 U1783 ( .A1(n6917), .A2(\mem[110][8] ), .B1(n6966), .B2(
        \mem[114][8] ), .ZN(n5607) );
  AOI22D0 U1784 ( .A1(n6892), .A2(\mem[108][8] ), .B1(n6923), .B2(\mem[98][8] ), .ZN(n5606) );
  ND4D0 U1785 ( .A1(n5609), .A2(n5608), .A3(n5607), .A4(n5606), .ZN(n5620) );
  AOI22D0 U1786 ( .A1(n6982), .A2(\mem[66][8] ), .B1(n6912), .B2(\mem[120][8] ), .ZN(n5613) );
  AOI22D0 U1787 ( .A1(n6890), .A2(\mem[100][8] ), .B1(n6791), .B2(\mem[96][8] ), .ZN(n5612) );
  AOI22D0 U1788 ( .A1(n6859), .A2(\mem[116][8] ), .B1(n6935), .B2(
        \mem[127][8] ), .ZN(n5610) );
  ND4D0 U1789 ( .A1(n5613), .A2(n5612), .A3(n5611), .A4(n5610), .ZN(n5619) );
  AOI22D0 U1790 ( .A1(n6981), .A2(\mem[124][8] ), .B1(n6968), .B2(
        \mem[105][8] ), .ZN(n5617) );
  AOI22D0 U1791 ( .A1(n6991), .A2(\mem[84][8] ), .B1(n6847), .B2(\mem[89][8] ), 
        .ZN(n5616) );
  AOI22D0 U1792 ( .A1(n6983), .A2(\mem[112][8] ), .B1(n6992), .B2(
        \mem[118][8] ), .ZN(n5615) );
  AOI22D0 U1793 ( .A1(n6905), .A2(\mem[123][8] ), .B1(n6542), .B2(\mem[82][8] ), .ZN(n5614) );
  ND4D0 U1794 ( .A1(n5617), .A2(n5616), .A3(n5615), .A4(n5614), .ZN(n5618) );
  NR4D0 U1795 ( .A1(n5621), .A2(n5620), .A3(n5619), .A4(n5618), .ZN(n5643) );
  AOI22D0 U1796 ( .A1(n6934), .A2(\mem[88][8] ), .B1(n6933), .B2(\mem[97][8] ), 
        .ZN(n5625) );
  AOI22D0 U1797 ( .A1(n6959), .A2(\mem[67][8] ), .B1(n6990), .B2(\mem[76][8] ), 
        .ZN(n5624) );
  AOI22D0 U1798 ( .A1(n6860), .A2(\mem[99][8] ), .B1(n6965), .B2(\mem[77][8] ), 
        .ZN(n5623) );
  AOI22D0 U1799 ( .A1(n6957), .A2(\mem[121][8] ), .B1(n6956), .B2(
        \mem[104][8] ), .ZN(n5622) );
  AOI22D0 U1800 ( .A1(n6809), .A2(\mem[73][8] ), .B1(n6993), .B2(\mem[117][8] ), .ZN(n5629) );
  AOI22D0 U1801 ( .A1(n6891), .A2(\mem[90][8] ), .B1(n6936), .B2(\mem[81][8] ), 
        .ZN(n5628) );
  AOI22D0 U1802 ( .A1(n6814), .A2(\mem[65][8] ), .B1(n6914), .B2(\mem[69][8] ), 
        .ZN(n5627) );
  AOI22D0 U1803 ( .A1(n6971), .A2(\mem[102][8] ), .B1(n6789), .B2(
        \mem[126][8] ), .ZN(n5626) );
  ND4D0 U1804 ( .A1(n5629), .A2(n5628), .A3(n5627), .A4(n5626), .ZN(n5640) );
  AOI22D0 U1805 ( .A1(n6989), .A2(\mem[70][8] ), .B1(n6879), .B2(\mem[122][8] ), .ZN(n5633) );
  AOI22D0 U1806 ( .A1(n6639), .A2(\mem[103][8] ), .B1(n6978), .B2(\mem[72][8] ), .ZN(n5631) );
  AOI22D0 U1807 ( .A1(n6928), .A2(\mem[71][8] ), .B1(n6925), .B2(\mem[109][8] ), .ZN(n5630) );
  ND4D0 U1808 ( .A1(n5633), .A2(n5632), .A3(n5631), .A4(n5630), .ZN(n5639) );
  AOI22D0 U1809 ( .A1(n6861), .A2(\mem[68][8] ), .B1(n6837), .B2(\mem[79][8] ), 
        .ZN(n5637) );
  AOI22D0 U1810 ( .A1(n6874), .A2(\mem[106][8] ), .B1(n6836), .B2(\mem[74][8] ), .ZN(n5636) );
  AOI22D0 U1811 ( .A1(n6448), .A2(\mem[64][8] ), .B1(n6873), .B2(\mem[94][8] ), 
        .ZN(n5635) );
  AOI22D0 U1812 ( .A1(n6868), .A2(\mem[107][8] ), .B1(n6869), .B2(
        \mem[113][8] ), .ZN(n5634) );
  ND4D0 U1813 ( .A1(n5637), .A2(n5636), .A3(n5635), .A4(n5634), .ZN(n5638) );
  NR4D0 U1814 ( .A1(n5641), .A2(n5640), .A3(n5639), .A4(n5638), .ZN(n5642) );
  AOI21D0 U1815 ( .A1(n5643), .A2(n5642), .B(n7004), .ZN(n5644) );
  AOI211D0 U1816 ( .A1(n6951), .A2(n5646), .B(n5645), .C(n5644), .ZN(n5668) );
  AOI22D0 U1817 ( .A1(n6727), .A2(\mem[42][8] ), .B1(n6978), .B2(\mem[8][8] ), 
        .ZN(n5650) );
  AOI22D0 U1818 ( .A1(n6905), .A2(\mem[59][8] ), .B1(n6879), .B2(\mem[58][8] ), 
        .ZN(n5649) );
  AOI22D0 U1819 ( .A1(n6860), .A2(\mem[35][8] ), .B1(n6965), .B2(\mem[13][8] ), 
        .ZN(n5648) );
  AOI22D0 U1820 ( .A1(n6959), .A2(\mem[3][8] ), .B1(n6892), .B2(\mem[44][8] ), 
        .ZN(n5647) );
  ND4D0 U1821 ( .A1(n5650), .A2(n5649), .A3(n5648), .A4(n5647), .ZN(n5666) );
  AOI22D0 U1822 ( .A1(n6790), .A2(\mem[27][8] ), .B1(n6837), .B2(\mem[15][8] ), 
        .ZN(n5654) );
  AOI22D0 U1823 ( .A1(n6748), .A2(\mem[41][8] ), .B1(n6990), .B2(\mem[12][8] ), 
        .ZN(n5653) );
  AOI22D0 U1824 ( .A1(n6953), .A2(\mem[47][8] ), .B1(n6992), .B2(\mem[54][8] ), 
        .ZN(n5652) );
  AOI22D0 U1825 ( .A1(n6883), .A2(\mem[48][8] ), .B1(n6967), .B2(\mem[39][8] ), 
        .ZN(n5651) );
  ND4D0 U1826 ( .A1(n5654), .A2(n5653), .A3(n5652), .A4(n5651), .ZN(n5665) );
  AOI22D0 U1827 ( .A1(n6835), .A2(\mem[4][8] ), .B1(n6958), .B2(\mem[17][8] ), 
        .ZN(n5657) );
  AOI22D0 U1828 ( .A1(n6989), .A2(\mem[6][8] ), .B1(n6296), .B2(\mem[29][8] ), 
        .ZN(n5656) );
  AOI22D0 U1829 ( .A1(n6976), .A2(\mem[34][8] ), .B1(n6935), .B2(\mem[63][8] ), 
        .ZN(n5655) );
  AOI22D0 U1830 ( .A1(n6890), .A2(\mem[36][8] ), .B1(n6869), .B2(\mem[49][8] ), 
        .ZN(n5662) );
  AOI22D0 U1831 ( .A1(n6754), .A2(\mem[5][8] ), .B1(n6955), .B2(\mem[21][8] ), 
        .ZN(n5661) );
  AOI22D0 U1832 ( .A1(n6981), .A2(\mem[60][8] ), .B1(n6903), .B2(\mem[51][8] ), 
        .ZN(n5660) );
  AOI22D0 U1833 ( .A1(n6614), .A2(\mem[22][8] ), .B1(n6966), .B2(\mem[50][8] ), 
        .ZN(n5659) );
  ND4D0 U1834 ( .A1(n5662), .A2(n5661), .A3(n5660), .A4(n5659), .ZN(n5663) );
  NR4D0 U1835 ( .A1(n5666), .A2(n5665), .A3(n5664), .A4(n5663), .ZN(n5667) );
  AOI32D0 U1836 ( .A1(n5669), .A2(n5668), .A3(n5667), .B1(n6856), .B2(n5668), 
        .ZN(dout[8]) );
  AOI22D0 U1837 ( .A1(n6880), .A2(\mem[75][10] ), .B1(n6862), .B2(
        \mem[104][10] ), .ZN(n5673) );
  AOI22D0 U1838 ( .A1(n6835), .A2(\mem[68][10] ), .B1(n6913), .B2(
        \mem[91][10] ), .ZN(n5672) );
  AOI22D0 U1839 ( .A1(n6957), .A2(\mem[121][10] ), .B1(n6915), .B2(
        \mem[77][10] ), .ZN(n5671) );
  AOI22D0 U1840 ( .A1(n6830), .A2(\mem[71][10] ), .B1(n6814), .B2(
        \mem[65][10] ), .ZN(n5670) );
  ND4D0 U1841 ( .A1(n5673), .A2(n5672), .A3(n5671), .A4(n5670), .ZN(n5689) );
  AOI22D0 U1842 ( .A1(n6979), .A2(\mem[78][10] ), .B1(n6542), .B2(
        \mem[82][10] ), .ZN(n5677) );
  AOI22D0 U1843 ( .A1(n6773), .A2(\mem[100][10] ), .B1(n6925), .B2(
        \mem[109][10] ), .ZN(n5676) );
  AOI22D0 U1844 ( .A1(n6803), .A2(\mem[119][10] ), .B1(n6754), .B2(
        \mem[69][10] ), .ZN(n5675) );
  AOI22D0 U1845 ( .A1(n6802), .A2(\mem[88][10] ), .B1(n6774), .B2(
        \mem[113][10] ), .ZN(n5674) );
  AOI22D0 U1846 ( .A1(n6819), .A2(\mem[125][10] ), .B1(n6906), .B2(
        \mem[76][10] ), .ZN(n5681) );
  AOI22D0 U1847 ( .A1(n6872), .A2(\mem[70][10] ), .B1(n6916), .B2(
        \mem[85][10] ), .ZN(n5680) );
  AOI22D0 U1848 ( .A1(n6903), .A2(\mem[115][10] ), .B1(n6882), .B2(
        \mem[79][10] ), .ZN(n5679) );
  AOI22D0 U1849 ( .A1(n6859), .A2(\mem[116][10] ), .B1(n6804), .B2(
        \mem[83][10] ), .ZN(n5678) );
  ND4D0 U1850 ( .A1(n5681), .A2(n5680), .A3(n5679), .A4(n5678), .ZN(n5687) );
  AOI22D0 U1851 ( .A1(n6977), .A2(\mem[97][10] ), .B1(n6879), .B2(
        \mem[122][10] ), .ZN(n5685) );
  AOI22D0 U1852 ( .A1(n6530), .A2(\mem[123][10] ), .B1(n6995), .B2(
        \mem[87][10] ), .ZN(n5684) );
  AOI22D0 U1853 ( .A1(n6981), .A2(\mem[124][10] ), .B1(n6874), .B2(
        \mem[106][10] ), .ZN(n5682) );
  ND4D0 U1854 ( .A1(n5685), .A2(n5684), .A3(n5683), .A4(n5682), .ZN(n5686) );
  NR4D0 U1855 ( .A1(n5689), .A2(n5688), .A3(n5687), .A4(n5686), .ZN(n5841) );
  AOI22D0 U1856 ( .A1(n6775), .A2(\mem[172][10] ), .B1(n6860), .B2(
        \mem[163][10] ), .ZN(n5693) );
  AOI22D0 U1857 ( .A1(n6934), .A2(\mem[152][10] ), .B1(n6923), .B2(
        \mem[162][10] ), .ZN(n5692) );
  AOI22D0 U1858 ( .A1(n6970), .A2(\mem[144][10] ), .B1(n6913), .B2(
        \mem[155][10] ), .ZN(n5690) );
  ND4D0 U1859 ( .A1(n5693), .A2(n5692), .A3(n5691), .A4(n5690), .ZN(n5709) );
  AOI22D0 U1860 ( .A1(n6914), .A2(\mem[133][10] ), .B1(n6862), .B2(
        \mem[168][10] ), .ZN(n5697) );
  AOI22D0 U1861 ( .A1(n6868), .A2(\mem[171][10] ), .B1(n6922), .B2(
        \mem[157][10] ), .ZN(n5696) );
  AOI22D0 U1862 ( .A1(n6680), .A2(\mem[159][10] ), .B1(n6871), .B2(
        \mem[185][10] ), .ZN(n5695) );
  AOI22D0 U1863 ( .A1(n6883), .A2(\mem[176][10] ), .B1(n6966), .B2(
        \mem[178][10] ), .ZN(n5694) );
  ND4D0 U1864 ( .A1(n5697), .A2(n5696), .A3(n5695), .A4(n5694), .ZN(n5708) );
  AOI22D0 U1865 ( .A1(n6830), .A2(\mem[135][10] ), .B1(n6873), .B2(
        \mem[158][10] ), .ZN(n5701) );
  AOI22D0 U1866 ( .A1(n6952), .A2(\mem[150][10] ), .B1(n6958), .B2(
        \mem[145][10] ), .ZN(n5700) );
  AOI22D0 U1867 ( .A1(n6907), .A2(\mem[131][10] ), .B1(n6955), .B2(
        \mem[149][10] ), .ZN(n5699) );
  AOI22D0 U1868 ( .A1(n6953), .A2(\mem[175][10] ), .B1(n6889), .B2(
        \mem[156][10] ), .ZN(n5698) );
  AOI22D0 U1869 ( .A1(n6773), .A2(\mem[164][10] ), .B1(n6965), .B2(
        \mem[141][10] ), .ZN(n5705) );
  AOI22D0 U1870 ( .A1(n6933), .A2(\mem[161][10] ), .B1(n6542), .B2(
        \mem[146][10] ), .ZN(n5704) );
  AOI22D0 U1871 ( .A1(n6803), .A2(\mem[183][10] ), .B1(n6836), .B2(
        \mem[138][10] ), .ZN(n5703) );
  AOI22D0 U1872 ( .A1(n6891), .A2(\mem[154][10] ), .B1(n6809), .B2(
        \mem[137][10] ), .ZN(n5702) );
  ND4D0 U1873 ( .A1(n5705), .A2(n5704), .A3(n5703), .A4(n5702), .ZN(n5706) );
  NR4D0 U1874 ( .A1(n5709), .A2(n5708), .A3(n5707), .A4(n5706), .ZN(n5731) );
  AOI22D0 U1875 ( .A1(n6747), .A2(\mem[148][10] ), .B1(n6912), .B2(
        \mem[184][10] ), .ZN(n5713) );
  AOI22D0 U1876 ( .A1(n6870), .A2(\mem[188][10] ), .B1(n6733), .B2(
        \mem[186][10] ), .ZN(n5711) );
  AOI22D0 U1877 ( .A1(n6905), .A2(\mem[187][10] ), .B1(n6760), .B2(
        \mem[173][10] ), .ZN(n5710) );
  ND4D0 U1878 ( .A1(n5713), .A2(n5712), .A3(n5711), .A4(n5710), .ZN(n5729) );
  AOI22D0 U1879 ( .A1(n6917), .A2(\mem[174][10] ), .B1(n6926), .B2(
        \mem[129][10] ), .ZN(n5717) );
  AOI22D0 U1880 ( .A1(n6967), .A2(\mem[167][10] ), .B1(n6738), .B2(
        \mem[165][10] ), .ZN(n5716) );
  AOI22D0 U1881 ( .A1(n6835), .A2(\mem[132][10] ), .B1(n6874), .B2(
        \mem[170][10] ), .ZN(n5715) );
  AOI22D0 U1882 ( .A1(n6979), .A2(\mem[142][10] ), .B1(n6992), .B2(
        \mem[182][10] ), .ZN(n5714) );
  ND4D0 U1883 ( .A1(n5717), .A2(n5716), .A3(n5715), .A4(n5714), .ZN(n5728) );
  AOI22D0 U1884 ( .A1(n6847), .A2(\mem[153][10] ), .B1(n6748), .B2(
        \mem[169][10] ), .ZN(n5721) );
  AOI22D0 U1885 ( .A1(n6888), .A2(\mem[128][10] ), .B1(n6491), .B2(
        \mem[179][10] ), .ZN(n5720) );
  AOI22D0 U1886 ( .A1(n6872), .A2(\mem[134][10] ), .B1(n6994), .B2(
        \mem[190][10] ), .ZN(n5719) );
  AOI22D0 U1887 ( .A1(n6880), .A2(\mem[139][10] ), .B1(n6728), .B2(
        \mem[180][10] ), .ZN(n5718) );
  ND4D0 U1888 ( .A1(n5721), .A2(n5720), .A3(n5719), .A4(n5718), .ZN(n5727) );
  AOI22D0 U1889 ( .A1(n6982), .A2(\mem[130][10] ), .B1(n6906), .B2(
        \mem[140][10] ), .ZN(n5725) );
  AOI22D0 U1890 ( .A1(n6995), .A2(\mem[151][10] ), .B1(n6935), .B2(
        \mem[191][10] ), .ZN(n5724) );
  AOI22D0 U1891 ( .A1(n6819), .A2(\mem[189][10] ), .B1(n6563), .B2(
        \mem[136][10] ), .ZN(n5723) );
  AOI22D0 U1892 ( .A1(n6659), .A2(\mem[181][10] ), .B1(n6774), .B2(
        \mem[177][10] ), .ZN(n5722) );
  ND4D0 U1893 ( .A1(n5725), .A2(n5724), .A3(n5723), .A4(n5722), .ZN(n5726) );
  NR4D0 U1894 ( .A1(n5729), .A2(n5728), .A3(n5727), .A4(n5726), .ZN(n5730) );
  CKND2D0 U1895 ( .A1(n5731), .A2(n5730), .ZN(n5818) );
  AOI22D0 U1896 ( .A1(n6814), .A2(\mem[1][10] ), .B1(n6988), .B2(\mem[63][10] ), .ZN(n5734) );
  AOI22D0 U1897 ( .A1(n6830), .A2(\mem[7][10] ), .B1(n6959), .B2(\mem[3][10] ), 
        .ZN(n5733) );
  AOI22D0 U1898 ( .A1(n6924), .A2(\mem[32][10] ), .B1(n6964), .B2(
        \mem[30][10] ), .ZN(n5732) );
  ND4D0 U1899 ( .A1(n5735), .A2(n5734), .A3(n5733), .A4(n5732), .ZN(n5751) );
  AOI22D0 U1900 ( .A1(n6922), .A2(\mem[29][10] ), .B1(n6728), .B2(
        \mem[52][10] ), .ZN(n5739) );
  AOI22D0 U1901 ( .A1(n6530), .A2(\mem[59][10] ), .B1(n6698), .B2(\mem[2][10] ), .ZN(n5738) );
  AOI22D0 U1902 ( .A1(n6903), .A2(\mem[51][10] ), .B1(n6658), .B2(
        \mem[50][10] ), .ZN(n5737) );
  AOI22D0 U1903 ( .A1(n6773), .A2(\mem[36][10] ), .B1(n6868), .B2(
        \mem[43][10] ), .ZN(n5736) );
  ND4D0 U1904 ( .A1(n5739), .A2(n5738), .A3(n5737), .A4(n5736), .ZN(n5750) );
  AOI22D0 U1905 ( .A1(n6879), .A2(\mem[58][10] ), .B1(n6915), .B2(
        \mem[13][10] ), .ZN(n5743) );
  AOI22D0 U1906 ( .A1(n6970), .A2(\mem[16][10] ), .B1(n6906), .B2(
        \mem[12][10] ), .ZN(n5742) );
  AOI22D0 U1907 ( .A1(n6179), .A2(\mem[47][10] ), .B1(n6880), .B2(
        \mem[11][10] ), .ZN(n5741) );
  AOI22D0 U1908 ( .A1(n6165), .A2(\mem[46][10] ), .B1(n6933), .B2(
        \mem[33][10] ), .ZN(n5740) );
  ND4D0 U1909 ( .A1(n5743), .A2(n5742), .A3(n5741), .A4(n5740), .ZN(n5749) );
  AOI22D0 U1910 ( .A1(n6981), .A2(\mem[60][10] ), .B1(n6835), .B2(\mem[4][10] ), .ZN(n5747) );
  AOI22D0 U1911 ( .A1(n6819), .A2(\mem[61][10] ), .B1(n6993), .B2(
        \mem[53][10] ), .ZN(n5746) );
  AOI22D0 U1912 ( .A1(n6952), .A2(\mem[22][10] ), .B1(n6784), .B2(
        \mem[28][10] ), .ZN(n5745) );
  ND4D0 U1913 ( .A1(n5747), .A2(n5746), .A3(n5745), .A4(n5744), .ZN(n5748) );
  NR4D0 U1914 ( .A1(n5751), .A2(n5750), .A3(n5749), .A4(n5748), .ZN(n5773) );
  AOI22D0 U1915 ( .A1(n6891), .A2(\mem[26][10] ), .B1(n6862), .B2(
        \mem[40][10] ), .ZN(n5755) );
  AOI22D0 U1916 ( .A1(n6639), .A2(\mem[39][10] ), .B1(n6727), .B2(
        \mem[42][10] ), .ZN(n5754) );
  AOI22D0 U1917 ( .A1(n6957), .A2(\mem[57][10] ), .B1(n6760), .B2(
        \mem[45][10] ), .ZN(n5753) );
  AOI22D0 U1918 ( .A1(n6901), .A2(\mem[9][10] ), .B1(n6738), .B2(\mem[37][10] ), .ZN(n5752) );
  ND4D0 U1919 ( .A1(n5755), .A2(n5754), .A3(n5753), .A4(n5752), .ZN(n5771) );
  AOI22D0 U1920 ( .A1(n6872), .A2(\mem[6][10] ), .B1(n6983), .B2(\mem[48][10] ), .ZN(n5759) );
  AOI22D0 U1921 ( .A1(n6847), .A2(\mem[25][10] ), .B1(n6954), .B2(
        \mem[10][10] ), .ZN(n5758) );
  AOI22D0 U1922 ( .A1(n6802), .A2(\mem[24][10] ), .B1(n6863), .B2(
        \mem[55][10] ), .ZN(n5757) );
  AOI22D0 U1923 ( .A1(n6971), .A2(\mem[38][10] ), .B1(n6774), .B2(
        \mem[49][10] ), .ZN(n5756) );
  ND4D0 U1924 ( .A1(n5759), .A2(n5758), .A3(n5757), .A4(n5756), .ZN(n5770) );
  AOI22D0 U1925 ( .A1(n6968), .A2(\mem[41][10] ), .B1(n6882), .B2(
        \mem[15][10] ), .ZN(n5763) );
  AOI22D0 U1926 ( .A1(n6914), .A2(\mem[5][10] ), .B1(n5966), .B2(\mem[31][10] ), .ZN(n5762) );
  AOI22D0 U1927 ( .A1(n6888), .A2(\mem[0][10] ), .B1(n6936), .B2(\mem[17][10] ), .ZN(n5761) );
  AOI22D0 U1928 ( .A1(n6969), .A2(\mem[18][10] ), .B1(n6904), .B2(
        \mem[19][10] ), .ZN(n5760) );
  ND4D0 U1929 ( .A1(n5763), .A2(n5762), .A3(n5761), .A4(n5760), .ZN(n5769) );
  AOI22D0 U1930 ( .A1(n6913), .A2(\mem[27][10] ), .B1(n6707), .B2(
        \mem[23][10] ), .ZN(n5767) );
  AOI22D0 U1931 ( .A1(n6979), .A2(\mem[14][10] ), .B1(n6828), .B2(
        \mem[56][10] ), .ZN(n5766) );
  AOI22D0 U1932 ( .A1(n6978), .A2(\mem[8][10] ), .B1(n6174), .B2(\mem[54][10] ), .ZN(n5764) );
  ND4D0 U1933 ( .A1(n5767), .A2(n5766), .A3(n5765), .A4(n5764), .ZN(n5768) );
  NR4D0 U1934 ( .A1(n5771), .A2(n5770), .A3(n5769), .A4(n5768), .ZN(n5772) );
  AOI21D0 U1935 ( .A1(n5773), .A2(n5772), .B(n6856), .ZN(n5817) );
  AOI22D0 U1936 ( .A1(n6803), .A2(\mem[247][10] ), .B1(n6754), .B2(
        \mem[197][10] ), .ZN(n5777) );
  AOI22D0 U1937 ( .A1(n6542), .A2(\mem[210][10] ), .B1(n6906), .B2(
        \mem[204][10] ), .ZN(n5776) );
  AOI22D0 U1938 ( .A1(n6991), .A2(\mem[212][10] ), .B1(n6491), .B2(
        \mem[243][10] ), .ZN(n5775) );
  AOI22D0 U1939 ( .A1(n6967), .A2(\mem[231][10] ), .B1(n6922), .B2(
        \mem[221][10] ), .ZN(n5774) );
  ND4D0 U1940 ( .A1(n5777), .A2(n5776), .A3(n5775), .A4(n5774), .ZN(n5793) );
  AOI22D0 U1941 ( .A1(n6835), .A2(\mem[196][10] ), .B1(n6968), .B2(
        \mem[233][10] ), .ZN(n5781) );
  AOI22D0 U1942 ( .A1(n6775), .A2(\mem[236][10] ), .B1(n6905), .B2(
        \mem[251][10] ), .ZN(n5780) );
  AOI22D0 U1943 ( .A1(n6525), .A2(\mem[227][10] ), .B1(n6955), .B2(
        \mem[213][10] ), .ZN(n5779) );
  AOI22D0 U1944 ( .A1(n6830), .A2(\mem[199][10] ), .B1(n6959), .B2(
        \mem[195][10] ), .ZN(n5778) );
  AOI22D0 U1945 ( .A1(n6760), .A2(\mem[237][10] ), .B1(n6978), .B2(
        \mem[200][10] ), .ZN(n5785) );
  AOI22D0 U1946 ( .A1(n6680), .A2(\mem[223][10] ), .B1(n6988), .B2(
        \mem[255][10] ), .ZN(n5784) );
  AOI22D0 U1947 ( .A1(n6165), .A2(\mem[238][10] ), .B1(n6842), .B2(
        \mem[218][10] ), .ZN(n5783) );
  AOI22D0 U1948 ( .A1(n6970), .A2(\mem[208][10] ), .B1(n6954), .B2(
        \mem[202][10] ), .ZN(n5782) );
  ND4D0 U1949 ( .A1(n5785), .A2(n5784), .A3(n5783), .A4(n5782), .ZN(n5791) );
  AOI22D0 U1950 ( .A1(n6773), .A2(\mem[228][10] ), .B1(n6727), .B2(
        \mem[234][10] ), .ZN(n5789) );
  AOI22D0 U1951 ( .A1(n6880), .A2(\mem[203][10] ), .B1(n6989), .B2(
        \mem[198][10] ), .ZN(n5787) );
  AOI22D0 U1952 ( .A1(n6913), .A2(\mem[219][10] ), .B1(n6995), .B2(
        \mem[215][10] ), .ZN(n5786) );
  ND4D0 U1953 ( .A1(n5789), .A2(n5788), .A3(n5787), .A4(n5786), .ZN(n5790) );
  NR4D0 U1954 ( .A1(n5793), .A2(n5792), .A3(n5791), .A4(n5790), .ZN(n5815) );
  AOI22D0 U1955 ( .A1(n6847), .A2(\mem[217][10] ), .B1(n6828), .B2(
        \mem[248][10] ), .ZN(n5797) );
  AOI22D0 U1956 ( .A1(n6952), .A2(\mem[214][10] ), .B1(n6926), .B2(
        \mem[193][10] ), .ZN(n5796) );
  AOI22D0 U1957 ( .A1(n6784), .A2(\mem[220][10] ), .B1(n6983), .B2(
        \mem[240][10] ), .ZN(n5795) );
  AOI22D0 U1958 ( .A1(n6819), .A2(\mem[253][10] ), .B1(n6933), .B2(
        \mem[225][10] ), .ZN(n5794) );
  ND4D0 U1959 ( .A1(n5797), .A2(n5796), .A3(n5795), .A4(n5794), .ZN(n5813) );
  AOI22D0 U1960 ( .A1(n6870), .A2(\mem[252][10] ), .B1(n6804), .B2(
        \mem[211][10] ), .ZN(n5801) );
  AOI22D0 U1961 ( .A1(n6879), .A2(\mem[250][10] ), .B1(n6982), .B2(
        \mem[194][10] ), .ZN(n5800) );
  AOI22D0 U1962 ( .A1(n6448), .A2(\mem[192][10] ), .B1(n6924), .B2(
        \mem[224][10] ), .ZN(n5799) );
  AOI22D0 U1963 ( .A1(n6957), .A2(\mem[249][10] ), .B1(n6774), .B2(
        \mem[241][10] ), .ZN(n5798) );
  ND4D0 U1964 ( .A1(n5801), .A2(n5800), .A3(n5799), .A4(n5798), .ZN(n5812) );
  AOI22D0 U1965 ( .A1(n6789), .A2(\mem[254][10] ), .B1(n6738), .B2(
        \mem[229][10] ), .ZN(n5805) );
  AOI22D0 U1966 ( .A1(n6179), .A2(\mem[239][10] ), .B1(n6964), .B2(
        \mem[222][10] ), .ZN(n5804) );
  AOI22D0 U1967 ( .A1(n6868), .A2(\mem[235][10] ), .B1(n6882), .B2(
        \mem[207][10] ), .ZN(n5803) );
  AOI22D0 U1968 ( .A1(n6809), .A2(\mem[201][10] ), .B1(n6174), .B2(
        \mem[246][10] ), .ZN(n5802) );
  ND4D0 U1969 ( .A1(n5805), .A2(n5804), .A3(n5803), .A4(n5802), .ZN(n5811) );
  AOI22D0 U1970 ( .A1(n6923), .A2(\mem[226][10] ), .B1(n6965), .B2(
        \mem[205][10] ), .ZN(n5808) );
  AOI22D0 U1971 ( .A1(n6829), .A2(\mem[230][10] ), .B1(n6956), .B2(
        \mem[232][10] ), .ZN(n5807) );
  AOI22D0 U1972 ( .A1(n6993), .A2(\mem[245][10] ), .B1(n6728), .B2(
        \mem[244][10] ), .ZN(n5806) );
  ND4D0 U1973 ( .A1(n5809), .A2(n5808), .A3(n5807), .A4(n5806), .ZN(n5810) );
  NR4D0 U1974 ( .A1(n5813), .A2(n5812), .A3(n5811), .A4(n5810), .ZN(n5814) );
  AOI21D0 U1975 ( .A1(n5815), .A2(n5814), .B(n6945), .ZN(n5816) );
  AOI211D0 U1976 ( .A1(n6951), .A2(n5818), .B(n5817), .C(n5816), .ZN(n5840) );
  AOI22D0 U1977 ( .A1(n6966), .A2(\mem[114][10] ), .B1(n6988), .B2(
        \mem[127][10] ), .ZN(n5822) );
  AOI22D0 U1978 ( .A1(n6847), .A2(\mem[89][10] ), .B1(n6828), .B2(
        \mem[120][10] ), .ZN(n5821) );
  AOI22D0 U1979 ( .A1(n6924), .A2(\mem[96][10] ), .B1(n6964), .B2(
        \mem[94][10] ), .ZN(n5820) );
  AOI22D0 U1980 ( .A1(n6836), .A2(\mem[74][10] ), .B1(n6738), .B2(
        \mem[101][10] ), .ZN(n5819) );
  ND4D0 U1981 ( .A1(n5822), .A2(n5821), .A3(n5820), .A4(n5819), .ZN(n5838) );
  AOI22D0 U1982 ( .A1(n6775), .A2(\mem[108][10] ), .B1(n6923), .B2(
        \mem[98][10] ), .ZN(n5826) );
  AOI22D0 U1983 ( .A1(n6970), .A2(\mem[80][10] ), .B1(n6968), .B2(
        \mem[105][10] ), .ZN(n5825) );
  AOI22D0 U1984 ( .A1(n6639), .A2(\mem[103][10] ), .B1(n6993), .B2(
        \mem[117][10] ), .ZN(n5824) );
  ND4D0 U1985 ( .A1(n5826), .A2(n5825), .A3(n5824), .A4(n5823), .ZN(n5837) );
  AOI22D0 U1986 ( .A1(n6868), .A2(\mem[107][10] ), .B1(n6994), .B2(
        \mem[126][10] ), .ZN(n5830) );
  AOI22D0 U1987 ( .A1(n6784), .A2(\mem[92][10] ), .B1(n6680), .B2(
        \mem[95][10] ), .ZN(n5829) );
  AOI22D0 U1988 ( .A1(n6917), .A2(\mem[110][10] ), .B1(n6842), .B2(
        \mem[90][10] ), .ZN(n5828) );
  AOI22D0 U1989 ( .A1(n6907), .A2(\mem[67][10] ), .B1(n6698), .B2(
        \mem[66][10] ), .ZN(n5827) );
  ND4D0 U1990 ( .A1(n5830), .A2(n5829), .A3(n5828), .A4(n5827), .ZN(n5836) );
  AOI22D0 U1991 ( .A1(n6888), .A2(\mem[64][10] ), .B1(n6936), .B2(
        \mem[81][10] ), .ZN(n5834) );
  AOI22D0 U1992 ( .A1(n6563), .A2(\mem[72][10] ), .B1(n6992), .B2(
        \mem[118][10] ), .ZN(n5833) );
  AOI22D0 U1993 ( .A1(n6953), .A2(\mem[111][10] ), .B1(n6983), .B2(
        \mem[112][10] ), .ZN(n5832) );
  AOI22D0 U1994 ( .A1(n6952), .A2(\mem[86][10] ), .B1(n6991), .B2(
        \mem[84][10] ), .ZN(n5831) );
  ND4D0 U1995 ( .A1(n5834), .A2(n5833), .A3(n5832), .A4(n5831), .ZN(n5835) );
  NR4D0 U1996 ( .A1(n5838), .A2(n5837), .A3(n5836), .A4(n5835), .ZN(n5839) );
  AOI32D0 U1997 ( .A1(n5841), .A2(n5840), .A3(n5839), .B1(n7004), .B2(n5840), 
        .ZN(dout[10]) );
  AOI22D0 U1998 ( .A1(n6804), .A2(\mem[147][9] ), .B1(n6964), .B2(
        \mem[158][9] ), .ZN(n5845) );
  AOI22D0 U1999 ( .A1(n6525), .A2(\mem[163][9] ), .B1(n6847), .B2(
        \mem[153][9] ), .ZN(n5844) );
  AOI22D0 U2000 ( .A1(n6814), .A2(\mem[129][9] ), .B1(n6861), .B2(
        \mem[132][9] ), .ZN(n5843) );
  AOI22D0 U2001 ( .A1(n6773), .A2(\mem[164][9] ), .B1(n6789), .B2(
        \mem[190][9] ), .ZN(n5842) );
  ND4D0 U2002 ( .A1(n5845), .A2(n5844), .A3(n5843), .A4(n5842), .ZN(n5861) );
  AOI22D0 U2003 ( .A1(n6956), .A2(\mem[168][9] ), .B1(n6828), .B2(
        \mem[184][9] ), .ZN(n5849) );
  AOI22D0 U2004 ( .A1(n6892), .A2(\mem[172][9] ), .B1(n6967), .B2(
        \mem[167][9] ), .ZN(n5848) );
  AOI22D0 U2005 ( .A1(n6872), .A2(\mem[134][9] ), .B1(n6784), .B2(
        \mem[156][9] ), .ZN(n5847) );
  ND4D0 U2006 ( .A1(n5849), .A2(n5848), .A3(n5847), .A4(n5846), .ZN(n5860) );
  AOI22D0 U2007 ( .A1(n6954), .A2(\mem[138][9] ), .B1(n6882), .B2(
        \mem[143][9] ), .ZN(n5853) );
  AOI22D0 U2008 ( .A1(n6325), .A2(\mem[139][9] ), .B1(n6955), .B2(
        \mem[149][9] ), .ZN(n5852) );
  AOI22D0 U2009 ( .A1(n6803), .A2(\mem[183][9] ), .B1(n6871), .B2(
        \mem[185][9] ), .ZN(n5851) );
  AOI22D0 U2010 ( .A1(n6830), .A2(\mem[135][9] ), .B1(n6905), .B2(
        \mem[187][9] ), .ZN(n5850) );
  ND4D0 U2011 ( .A1(n5853), .A2(n5852), .A3(n5851), .A4(n5850), .ZN(n5859) );
  AOI22D0 U2012 ( .A1(n6952), .A2(\mem[150][9] ), .B1(n6988), .B2(
        \mem[191][9] ), .ZN(n5857) );
  AOI22D0 U2013 ( .A1(n6907), .A2(\mem[131][9] ), .B1(n6903), .B2(
        \mem[179][9] ), .ZN(n5856) );
  AOI22D0 U2014 ( .A1(n6977), .A2(\mem[161][9] ), .B1(n5966), .B2(
        \mem[159][9] ), .ZN(n5855) );
  AOI22D0 U2015 ( .A1(n6991), .A2(\mem[148][9] ), .B1(n6968), .B2(
        \mem[169][9] ), .ZN(n5854) );
  ND4D0 U2016 ( .A1(n5857), .A2(n5856), .A3(n5855), .A4(n5854), .ZN(n5858) );
  NR4D0 U2017 ( .A1(n5861), .A2(n5860), .A3(n5859), .A4(n5858), .ZN(n6014) );
  AOI22D0 U2018 ( .A1(n6977), .A2(\mem[97][9] ), .B1(n6982), .B2(\mem[66][9] ), 
        .ZN(n5865) );
  AOI22D0 U2019 ( .A1(n6952), .A2(\mem[86][9] ), .B1(n6760), .B2(\mem[109][9] ), .ZN(n5864) );
  AOI22D0 U2020 ( .A1(n6707), .A2(\mem[87][9] ), .B1(n6994), .B2(\mem[126][9] ), .ZN(n5863) );
  AOI22D0 U2021 ( .A1(n6928), .A2(\mem[71][9] ), .B1(n6965), .B2(\mem[77][9] ), 
        .ZN(n5862) );
  ND4D0 U2022 ( .A1(n5865), .A2(n5864), .A3(n5863), .A4(n5862), .ZN(n5881) );
  AOI22D0 U2023 ( .A1(n6790), .A2(\mem[91][9] ), .B1(n6954), .B2(\mem[74][9] ), 
        .ZN(n5869) );
  AOI22D0 U2024 ( .A1(n6802), .A2(\mem[88][9] ), .B1(n6926), .B2(\mem[65][9] ), 
        .ZN(n5868) );
  AOI22D0 U2025 ( .A1(n6861), .A2(\mem[68][9] ), .B1(n6891), .B2(\mem[90][9] ), 
        .ZN(n5867) );
  AOI22D0 U2026 ( .A1(n6988), .A2(\mem[127][9] ), .B1(n6862), .B2(
        \mem[104][9] ), .ZN(n5866) );
  ND4D0 U2027 ( .A1(n5869), .A2(n5868), .A3(n5867), .A4(n5866), .ZN(n5880) );
  AOI22D0 U2028 ( .A1(n6179), .A2(\mem[111][9] ), .B1(n6922), .B2(\mem[93][9] ), .ZN(n5872) );
  AOI22D0 U2029 ( .A1(n6658), .A2(\mem[114][9] ), .B1(n6828), .B2(
        \mem[120][9] ), .ZN(n5871) );
  AOI22D0 U2030 ( .A1(n6892), .A2(\mem[108][9] ), .B1(n6881), .B2(\mem[80][9] ), .ZN(n5870) );
  ND4D0 U2031 ( .A1(n5873), .A2(n5872), .A3(n5871), .A4(n5870), .ZN(n5879) );
  AOI22D0 U2032 ( .A1(n6784), .A2(\mem[92][9] ), .B1(n6774), .B2(\mem[113][9] ), .ZN(n5877) );
  AOI22D0 U2033 ( .A1(n6991), .A2(\mem[84][9] ), .B1(n5966), .B2(\mem[95][9] ), 
        .ZN(n5876) );
  AOI22D0 U2034 ( .A1(n6860), .A2(\mem[99][9] ), .B1(n6906), .B2(\mem[76][9] ), 
        .ZN(n5875) );
  AOI22D0 U2035 ( .A1(n6983), .A2(\mem[112][9] ), .B1(n6964), .B2(\mem[94][9] ), .ZN(n5874) );
  ND4D0 U2036 ( .A1(n5877), .A2(n5876), .A3(n5875), .A4(n5874), .ZN(n5878) );
  NR4D0 U2037 ( .A1(n5881), .A2(n5880), .A3(n5879), .A4(n5878), .ZN(n5903) );
  AOI22D0 U2038 ( .A1(n6880), .A2(\mem[75][9] ), .B1(n6791), .B2(\mem[96][9] ), 
        .ZN(n5885) );
  AOI22D0 U2039 ( .A1(n6773), .A2(\mem[100][9] ), .B1(n6809), .B2(\mem[73][9] ), .ZN(n5884) );
  AOI22D0 U2040 ( .A1(n6981), .A2(\mem[124][9] ), .B1(n6733), .B2(
        \mem[122][9] ), .ZN(n5883) );
  AOI22D0 U2041 ( .A1(n6904), .A2(\mem[83][9] ), .B1(n6978), .B2(\mem[72][9] ), 
        .ZN(n5882) );
  ND4D0 U2042 ( .A1(n5885), .A2(n5884), .A3(n5883), .A4(n5882), .ZN(n5901) );
  AOI22D0 U2043 ( .A1(n6868), .A2(\mem[107][9] ), .B1(n6993), .B2(
        \mem[117][9] ), .ZN(n5889) );
  AOI22D0 U2044 ( .A1(n6165), .A2(\mem[110][9] ), .B1(n6980), .B2(
        \mem[125][9] ), .ZN(n5888) );
  AOI22D0 U2045 ( .A1(n6989), .A2(\mem[70][9] ), .B1(n6888), .B2(\mem[64][9] ), 
        .ZN(n5887) );
  ND4D0 U2046 ( .A1(n5889), .A2(n5888), .A3(n5887), .A4(n5886), .ZN(n5900) );
  AOI22D0 U2047 ( .A1(n6905), .A2(\mem[123][9] ), .B1(n6491), .B2(
        \mem[115][9] ), .ZN(n5893) );
  AOI22D0 U2048 ( .A1(n6927), .A2(\mem[89][9] ), .B1(n6958), .B2(\mem[81][9] ), 
        .ZN(n5892) );
  AOI22D0 U2049 ( .A1(n6979), .A2(\mem[78][9] ), .B1(n6971), .B2(\mem[102][9] ), .ZN(n5891) );
  AOI22D0 U2050 ( .A1(n6639), .A2(\mem[103][9] ), .B1(n6727), .B2(
        \mem[106][9] ), .ZN(n5890) );
  ND4D0 U2051 ( .A1(n5893), .A2(n5892), .A3(n5891), .A4(n5890), .ZN(n5899) );
  AOI22D0 U2052 ( .A1(n6923), .A2(\mem[98][9] ), .B1(n6882), .B2(\mem[79][9] ), 
        .ZN(n5897) );
  AOI22D0 U2053 ( .A1(n6914), .A2(\mem[69][9] ), .B1(n6738), .B2(\mem[101][9] ), .ZN(n5896) );
  AOI22D0 U2054 ( .A1(n6907), .A2(\mem[67][9] ), .B1(n6957), .B2(\mem[121][9] ), .ZN(n5895) );
  AOI22D0 U2055 ( .A1(n6969), .A2(\mem[82][9] ), .B1(n6955), .B2(\mem[85][9] ), 
        .ZN(n5894) );
  ND4D0 U2056 ( .A1(n5897), .A2(n5896), .A3(n5895), .A4(n5894), .ZN(n5898) );
  NR4D0 U2057 ( .A1(n5901), .A2(n5900), .A3(n5899), .A4(n5898), .ZN(n5902) );
  CKND2D0 U2058 ( .A1(n5903), .A2(n5902), .ZN(n5991) );
  AOI22D0 U2059 ( .A1(n6842), .A2(\mem[26][9] ), .B1(n6809), .B2(\mem[9][9] ), 
        .ZN(n5907) );
  AOI22D0 U2060 ( .A1(n6977), .A2(\mem[33][9] ), .B1(n6754), .B2(\mem[5][9] ), 
        .ZN(n5906) );
  AOI22D0 U2061 ( .A1(n6789), .A2(\mem[62][9] ), .B1(n6774), .B2(\mem[49][9] ), 
        .ZN(n5905) );
  AOI22D0 U2062 ( .A1(n6892), .A2(\mem[44][9] ), .B1(n6982), .B2(\mem[2][9] ), 
        .ZN(n5904) );
  ND4D0 U2063 ( .A1(n5907), .A2(n5906), .A3(n5905), .A4(n5904), .ZN(n5923) );
  AOI22D0 U2064 ( .A1(n6979), .A2(\mem[14][9] ), .B1(n6880), .B2(\mem[11][9] ), 
        .ZN(n5911) );
  AOI22D0 U2065 ( .A1(n6917), .A2(\mem[46][9] ), .B1(n6995), .B2(\mem[23][9] ), 
        .ZN(n5910) );
  AOI22D0 U2066 ( .A1(n6905), .A2(\mem[59][9] ), .B1(n6913), .B2(\mem[27][9] ), 
        .ZN(n5908) );
  ND4D0 U2067 ( .A1(n5911), .A2(n5910), .A3(n5909), .A4(n5908), .ZN(n5922) );
  AOI22D0 U2068 ( .A1(n6819), .A2(\mem[61][9] ), .B1(n6983), .B2(\mem[48][9] ), 
        .ZN(n5915) );
  AOI22D0 U2069 ( .A1(n6953), .A2(\mem[47][9] ), .B1(n6903), .B2(\mem[51][9] ), 
        .ZN(n5914) );
  AOI22D0 U2070 ( .A1(n6874), .A2(\mem[42][9] ), .B1(n6904), .B2(\mem[19][9] ), 
        .ZN(n5913) );
  AOI22D0 U2071 ( .A1(n6680), .A2(\mem[31][9] ), .B1(n6916), .B2(\mem[21][9] ), 
        .ZN(n5912) );
  ND4D0 U2072 ( .A1(n5915), .A2(n5914), .A3(n5913), .A4(n5912), .ZN(n5921) );
  AOI22D0 U2073 ( .A1(n6907), .A2(\mem[3][9] ), .B1(n6971), .B2(\mem[38][9] ), 
        .ZN(n5919) );
  AOI22D0 U2074 ( .A1(n6728), .A2(\mem[52][9] ), .B1(n6992), .B2(\mem[54][9] ), 
        .ZN(n5918) );
  AOI22D0 U2075 ( .A1(n6993), .A2(\mem[53][9] ), .B1(n6924), .B2(\mem[32][9] ), 
        .ZN(n5917) );
  AOI22D0 U2076 ( .A1(n6296), .A2(\mem[29][9] ), .B1(n6968), .B2(\mem[41][9] ), 
        .ZN(n5916) );
  NR4D0 U2077 ( .A1(n5923), .A2(n5922), .A3(n5921), .A4(n5920), .ZN(n5945) );
  AOI22D0 U2078 ( .A1(n6934), .A2(\mem[24][9] ), .B1(n6868), .B2(\mem[43][9] ), 
        .ZN(n5927) );
  AOI22D0 U2079 ( .A1(n6870), .A2(\mem[60][9] ), .B1(n6836), .B2(\mem[10][9] ), 
        .ZN(n5926) );
  AOI22D0 U2080 ( .A1(n6614), .A2(\mem[22][9] ), .B1(n6814), .B2(\mem[1][9] ), 
        .ZN(n5925) );
  AOI22D0 U2081 ( .A1(n6860), .A2(\mem[35][9] ), .B1(n6733), .B2(\mem[58][9] ), 
        .ZN(n5924) );
  ND4D0 U2082 ( .A1(n5927), .A2(n5926), .A3(n5925), .A4(n5924), .ZN(n5943) );
  AOI22D0 U2083 ( .A1(n6658), .A2(\mem[50][9] ), .B1(n6738), .B2(\mem[37][9] ), 
        .ZN(n5931) );
  AOI22D0 U2084 ( .A1(n6989), .A2(\mem[6][9] ), .B1(n6760), .B2(\mem[45][9] ), 
        .ZN(n5929) );
  AOI22D0 U2085 ( .A1(n6862), .A2(\mem[40][9] ), .B1(n6906), .B2(\mem[12][9] ), 
        .ZN(n5928) );
  ND4D0 U2086 ( .A1(n5931), .A2(n5930), .A3(n5929), .A4(n5928), .ZN(n5942) );
  AOI22D0 U2087 ( .A1(n6861), .A2(\mem[4][9] ), .B1(n6871), .B2(\mem[57][9] ), 
        .ZN(n5935) );
  AOI22D0 U2088 ( .A1(n6936), .A2(\mem[17][9] ), .B1(n6965), .B2(\mem[13][9] ), 
        .ZN(n5934) );
  AOI22D0 U2089 ( .A1(n6928), .A2(\mem[7][9] ), .B1(n6828), .B2(\mem[56][9] ), 
        .ZN(n5933) );
  AOI22D0 U2090 ( .A1(n6888), .A2(\mem[0][9] ), .B1(n6863), .B2(\mem[55][9] ), 
        .ZN(n5932) );
  ND4D0 U2091 ( .A1(n5935), .A2(n5934), .A3(n5933), .A4(n5932), .ZN(n5941) );
  AOI22D0 U2092 ( .A1(n6991), .A2(\mem[20][9] ), .B1(n6978), .B2(\mem[8][9] ), 
        .ZN(n5939) );
  AOI22D0 U2093 ( .A1(n6969), .A2(\mem[18][9] ), .B1(n6964), .B2(\mem[30][9] ), 
        .ZN(n5938) );
  AOI22D0 U2094 ( .A1(n6773), .A2(\mem[36][9] ), .B1(n6882), .B2(\mem[15][9] ), 
        .ZN(n5937) );
  AOI22D0 U2095 ( .A1(n6881), .A2(\mem[16][9] ), .B1(n6988), .B2(\mem[63][9] ), 
        .ZN(n5936) );
  ND4D0 U2096 ( .A1(n5939), .A2(n5938), .A3(n5937), .A4(n5936), .ZN(n5940) );
  NR4D0 U2097 ( .A1(n5943), .A2(n5942), .A3(n5941), .A4(n5940), .ZN(n5944) );
  AOI21D0 U2098 ( .A1(n5945), .A2(n5944), .B(n6856), .ZN(n5990) );
  AOI22D0 U2099 ( .A1(n6542), .A2(\mem[210][9] ), .B1(n6970), .B2(
        \mem[208][9] ), .ZN(n5949) );
  AOI22D0 U2100 ( .A1(n6861), .A2(\mem[196][9] ), .B1(n6913), .B2(
        \mem[219][9] ), .ZN(n5948) );
  AOI22D0 U2101 ( .A1(n6891), .A2(\mem[218][9] ), .B1(n6982), .B2(
        \mem[194][9] ), .ZN(n5947) );
  AOI22D0 U2102 ( .A1(n6728), .A2(\mem[244][9] ), .B1(n6774), .B2(
        \mem[241][9] ), .ZN(n5946) );
  ND4D0 U2103 ( .A1(n5949), .A2(n5948), .A3(n5947), .A4(n5946), .ZN(n5965) );
  AOI22D0 U2104 ( .A1(n6979), .A2(\mem[206][9] ), .B1(n6954), .B2(
        \mem[202][9] ), .ZN(n5952) );
  AOI22D0 U2105 ( .A1(n6991), .A2(\mem[212][9] ), .B1(n6936), .B2(
        \mem[209][9] ), .ZN(n5951) );
  AOI22D0 U2106 ( .A1(n6993), .A2(\mem[245][9] ), .B1(n6748), .B2(
        \mem[233][9] ), .ZN(n5950) );
  ND4D0 U2107 ( .A1(n5953), .A2(n5952), .A3(n5951), .A4(n5950), .ZN(n5964) );
  AOI22D0 U2108 ( .A1(n6952), .A2(\mem[214][9] ), .B1(n6923), .B2(
        \mem[226][9] ), .ZN(n5957) );
  AOI22D0 U2109 ( .A1(n6905), .A2(\mem[251][9] ), .B1(n6933), .B2(
        \mem[225][9] ), .ZN(n5956) );
  AOI22D0 U2110 ( .A1(n6784), .A2(\mem[220][9] ), .B1(n6707), .B2(
        \mem[215][9] ), .ZN(n5955) );
  AOI22D0 U2111 ( .A1(n6957), .A2(\mem[249][9] ), .B1(n6882), .B2(
        \mem[207][9] ), .ZN(n5954) );
  ND4D0 U2112 ( .A1(n5957), .A2(n5956), .A3(n5955), .A4(n5954), .ZN(n5963) );
  AOI22D0 U2113 ( .A1(n6802), .A2(\mem[216][9] ), .B1(n6847), .B2(
        \mem[217][9] ), .ZN(n5961) );
  AOI22D0 U2114 ( .A1(n6863), .A2(\mem[247][9] ), .B1(n6903), .B2(
        \mem[243][9] ), .ZN(n5960) );
  AOI22D0 U2115 ( .A1(n6814), .A2(\mem[193][9] ), .B1(n6966), .B2(
        \mem[242][9] ), .ZN(n5959) );
  AOI22D0 U2116 ( .A1(n6917), .A2(\mem[238][9] ), .B1(n6789), .B2(
        \mem[254][9] ), .ZN(n5958) );
  ND4D0 U2117 ( .A1(n5961), .A2(n5960), .A3(n5959), .A4(n5958), .ZN(n5962) );
  NR4D0 U2118 ( .A1(n5965), .A2(n5964), .A3(n5963), .A4(n5962), .ZN(n5988) );
  AOI22D0 U2119 ( .A1(n6829), .A2(\mem[230][9] ), .B1(n6733), .B2(
        \mem[250][9] ), .ZN(n5970) );
  AOI22D0 U2120 ( .A1(n6860), .A2(\mem[227][9] ), .B1(n5966), .B2(
        \mem[223][9] ), .ZN(n5969) );
  AOI22D0 U2121 ( .A1(n6563), .A2(\mem[200][9] ), .B1(n6906), .B2(
        \mem[204][9] ), .ZN(n5968) );
  ND4D0 U2122 ( .A1(n5970), .A2(n5969), .A3(n5968), .A4(n5967), .ZN(n5986) );
  AOI22D0 U2123 ( .A1(n6989), .A2(\mem[198][9] ), .B1(n6809), .B2(
        \mem[201][9] ), .ZN(n5974) );
  AOI22D0 U2124 ( .A1(n6980), .A2(\mem[253][9] ), .B1(n6760), .B2(
        \mem[237][9] ), .ZN(n5973) );
  AOI22D0 U2125 ( .A1(n6981), .A2(\mem[252][9] ), .B1(n6988), .B2(
        \mem[255][9] ), .ZN(n5972) );
  AOI22D0 U2126 ( .A1(n6868), .A2(\mem[235][9] ), .B1(n6992), .B2(
        \mem[246][9] ), .ZN(n5971) );
  ND4D0 U2127 ( .A1(n5974), .A2(n5973), .A3(n5972), .A4(n5971), .ZN(n5985) );
  AOI22D0 U2128 ( .A1(n6914), .A2(\mem[197][9] ), .B1(n6904), .B2(
        \mem[211][9] ), .ZN(n5978) );
  AOI22D0 U2129 ( .A1(n6922), .A2(\mem[221][9] ), .B1(n6902), .B2(
        \mem[229][9] ), .ZN(n5977) );
  AOI22D0 U2130 ( .A1(n6892), .A2(\mem[236][9] ), .B1(n6964), .B2(
        \mem[222][9] ), .ZN(n5976) );
  AOI22D0 U2131 ( .A1(n6953), .A2(\mem[239][9] ), .B1(n6888), .B2(
        \mem[192][9] ), .ZN(n5975) );
  ND4D0 U2132 ( .A1(n5978), .A2(n5977), .A3(n5976), .A4(n5975), .ZN(n5984) );
  AOI22D0 U2133 ( .A1(n6880), .A2(\mem[203][9] ), .B1(n6639), .B2(
        \mem[231][9] ), .ZN(n5982) );
  AOI22D0 U2134 ( .A1(n6874), .A2(\mem[234][9] ), .B1(n6965), .B2(
        \mem[205][9] ), .ZN(n5981) );
  AOI22D0 U2135 ( .A1(n6959), .A2(\mem[195][9] ), .B1(n6956), .B2(
        \mem[232][9] ), .ZN(n5980) );
  AOI22D0 U2136 ( .A1(n6916), .A2(\mem[213][9] ), .B1(n6828), .B2(
        \mem[248][9] ), .ZN(n5979) );
  ND4D0 U2137 ( .A1(n5982), .A2(n5981), .A3(n5980), .A4(n5979), .ZN(n5983) );
  NR4D0 U2138 ( .A1(n5986), .A2(n5985), .A3(n5984), .A4(n5983), .ZN(n5987) );
  AOI21D0 U2139 ( .A1(n5988), .A2(n5987), .B(n6945), .ZN(n5989) );
  AOI211D0 U2140 ( .A1(n6164), .A2(n5991), .B(n5990), .C(n5989), .ZN(n6013) );
  AOI22D0 U2141 ( .A1(n6993), .A2(\mem[181][9] ), .B1(n6958), .B2(
        \mem[145][9] ), .ZN(n5994) );
  AOI22D0 U2142 ( .A1(n6980), .A2(\mem[189][9] ), .B1(n6922), .B2(
        \mem[157][9] ), .ZN(n5993) );
  AOI22D0 U2143 ( .A1(n6728), .A2(\mem[180][9] ), .B1(n6902), .B2(
        \mem[165][9] ), .ZN(n5992) );
  ND4D0 U2144 ( .A1(n5995), .A2(n5994), .A3(n5993), .A4(n5992), .ZN(n6011) );
  AOI22D0 U2145 ( .A1(n6934), .A2(\mem[152][9] ), .B1(n6733), .B2(
        \mem[186][9] ), .ZN(n5999) );
  AOI22D0 U2146 ( .A1(n6870), .A2(\mem[188][9] ), .B1(n6978), .B2(
        \mem[136][9] ), .ZN(n5998) );
  AOI22D0 U2147 ( .A1(n6982), .A2(\mem[130][9] ), .B1(n6990), .B2(
        \mem[140][9] ), .ZN(n5997) );
  AOI22D0 U2148 ( .A1(n6965), .A2(\mem[141][9] ), .B1(n6760), .B2(
        \mem[173][9] ), .ZN(n5996) );
  ND4D0 U2149 ( .A1(n5999), .A2(n5998), .A3(n5997), .A4(n5996), .ZN(n6010) );
  AOI22D0 U2150 ( .A1(n6979), .A2(\mem[142][9] ), .B1(n6888), .B2(
        \mem[128][9] ), .ZN(n6003) );
  AOI22D0 U2151 ( .A1(n6953), .A2(\mem[175][9] ), .B1(n6874), .B2(
        \mem[170][9] ), .ZN(n6002) );
  AOI22D0 U2152 ( .A1(n6917), .A2(\mem[174][9] ), .B1(n6869), .B2(
        \mem[177][9] ), .ZN(n6001) );
  AOI22D0 U2153 ( .A1(n6971), .A2(\mem[166][9] ), .B1(n6970), .B2(
        \mem[144][9] ), .ZN(n6000) );
  ND4D0 U2154 ( .A1(n6003), .A2(n6002), .A3(n6001), .A4(n6000), .ZN(n6009) );
  AOI22D0 U2155 ( .A1(n6868), .A2(\mem[171][9] ), .B1(n6969), .B2(
        \mem[146][9] ), .ZN(n6007) );
  AOI22D0 U2156 ( .A1(n6809), .A2(\mem[137][9] ), .B1(n6992), .B2(
        \mem[182][9] ), .ZN(n6006) );
  AOI22D0 U2157 ( .A1(n6891), .A2(\mem[154][9] ), .B1(n6995), .B2(
        \mem[151][9] ), .ZN(n6005) );
  ND4D0 U2158 ( .A1(n6007), .A2(n6006), .A3(n6005), .A4(n6004), .ZN(n6008) );
  NR4D0 U2159 ( .A1(n6011), .A2(n6010), .A3(n6009), .A4(n6008), .ZN(n6012) );
  AOI32D0 U2160 ( .A1(n6014), .A2(n6013), .A3(n6012), .B1(n6188), .B2(n6013), 
        .ZN(dout[9]) );
  AOI22D0 U2161 ( .A1(n6890), .A2(\mem[164][6] ), .B1(n6979), .B2(
        \mem[142][6] ), .ZN(n6018) );
  AOI22D0 U2162 ( .A1(n6754), .A2(\mem[133][6] ), .B1(n6912), .B2(
        \mem[184][6] ), .ZN(n6017) );
  AOI22D0 U2163 ( .A1(n6614), .A2(\mem[150][6] ), .B1(n6964), .B2(
        \mem[158][6] ), .ZN(n6016) );
  AOI22D0 U2164 ( .A1(n6927), .A2(\mem[153][6] ), .B1(n6904), .B2(
        \mem[147][6] ), .ZN(n6015) );
  ND4D0 U2165 ( .A1(n6018), .A2(n6017), .A3(n6016), .A4(n6015), .ZN(n6034) );
  AOI22D0 U2166 ( .A1(n6957), .A2(\mem[185][6] ), .B1(n6882), .B2(
        \mem[143][6] ), .ZN(n6022) );
  AOI22D0 U2167 ( .A1(n6928), .A2(\mem[135][6] ), .B1(n6889), .B2(
        \mem[156][6] ), .ZN(n6021) );
  AOI22D0 U2168 ( .A1(n6658), .A2(\mem[178][6] ), .B1(n6748), .B2(
        \mem[169][6] ), .ZN(n6019) );
  ND4D0 U2169 ( .A1(n6022), .A2(n6021), .A3(n6020), .A4(n6019), .ZN(n6033) );
  AOI22D0 U2170 ( .A1(n6915), .A2(\mem[141][6] ), .B1(n6906), .B2(
        \mem[140][6] ), .ZN(n6026) );
  AOI22D0 U2171 ( .A1(n6881), .A2(\mem[144][6] ), .B1(n6888), .B2(
        \mem[128][6] ), .ZN(n6025) );
  AOI22D0 U2172 ( .A1(n6491), .A2(\mem[179][6] ), .B1(n6791), .B2(
        \mem[160][6] ), .ZN(n6024) );
  AOI22D0 U2173 ( .A1(n6728), .A2(\mem[180][6] ), .B1(n6869), .B2(
        \mem[177][6] ), .ZN(n6023) );
  ND4D0 U2174 ( .A1(n6026), .A2(n6025), .A3(n6024), .A4(n6023), .ZN(n6032) );
  AOI22D0 U2175 ( .A1(n6959), .A2(\mem[131][6] ), .B1(n6954), .B2(
        \mem[138][6] ), .ZN(n6030) );
  AOI22D0 U2176 ( .A1(n6989), .A2(\mem[134][6] ), .B1(n6902), .B2(
        \mem[165][6] ), .ZN(n6029) );
  AOI22D0 U2177 ( .A1(n6980), .A2(\mem[189][6] ), .B1(n6925), .B2(
        \mem[173][6] ), .ZN(n6028) );
  ND4D0 U2178 ( .A1(n6030), .A2(n6029), .A3(n6028), .A4(n6027), .ZN(n6031) );
  NR4D0 U2179 ( .A1(n6034), .A2(n6033), .A3(n6032), .A4(n6031), .ZN(n6191) );
  AOI22D0 U2180 ( .A1(n6179), .A2(\mem[111][6] ), .B1(n6905), .B2(
        \mem[123][6] ), .ZN(n6038) );
  AOI22D0 U2181 ( .A1(n6954), .A2(\mem[74][6] ), .B1(n6873), .B2(\mem[94][6] ), 
        .ZN(n6037) );
  AOI22D0 U2182 ( .A1(n6791), .A2(\mem[96][6] ), .B1(n6837), .B2(\mem[79][6] ), 
        .ZN(n6036) );
  AOI22D0 U2183 ( .A1(n6874), .A2(\mem[106][6] ), .B1(n6925), .B2(
        \mem[109][6] ), .ZN(n6035) );
  ND4D0 U2184 ( .A1(n6038), .A2(n6037), .A3(n6036), .A4(n6035), .ZN(n6054) );
  AOI22D0 U2185 ( .A1(n6983), .A2(\mem[112][6] ), .B1(n6728), .B2(
        \mem[116][6] ), .ZN(n6042) );
  AOI22D0 U2186 ( .A1(n6639), .A2(\mem[103][6] ), .B1(n6904), .B2(\mem[83][6] ), .ZN(n6041) );
  AOI22D0 U2187 ( .A1(n6928), .A2(\mem[71][6] ), .B1(n6889), .B2(\mem[92][6] ), 
        .ZN(n6040) );
  AOI22D0 U2188 ( .A1(n6802), .A2(\mem[88][6] ), .B1(n6868), .B2(\mem[107][6] ), .ZN(n6039) );
  ND4D0 U2189 ( .A1(n6042), .A2(n6041), .A3(n6040), .A4(n6039), .ZN(n6053) );
  AOI22D0 U2190 ( .A1(n6991), .A2(\mem[84][6] ), .B1(n6860), .B2(\mem[99][6] ), 
        .ZN(n6046) );
  AOI22D0 U2191 ( .A1(n6809), .A2(\mem[73][6] ), .B1(n6828), .B2(\mem[120][6] ), .ZN(n6045) );
  AOI22D0 U2192 ( .A1(n6903), .A2(\mem[115][6] ), .B1(n6174), .B2(
        \mem[118][6] ), .ZN(n6044) );
  ND4D0 U2193 ( .A1(n6046), .A2(n6045), .A3(n6044), .A4(n6043), .ZN(n6052) );
  AOI22D0 U2194 ( .A1(n6803), .A2(\mem[119][6] ), .B1(n6956), .B2(
        \mem[104][6] ), .ZN(n6050) );
  AOI22D0 U2195 ( .A1(n6789), .A2(\mem[126][6] ), .B1(n6748), .B2(
        \mem[105][6] ), .ZN(n6049) );
  AOI22D0 U2196 ( .A1(n6614), .A2(\mem[86][6] ), .B1(n6835), .B2(\mem[68][6] ), 
        .ZN(n6048) );
  AOI22D0 U2197 ( .A1(n6980), .A2(\mem[125][6] ), .B1(n6995), .B2(\mem[87][6] ), .ZN(n6047) );
  ND4D0 U2198 ( .A1(n6050), .A2(n6049), .A3(n6048), .A4(n6047), .ZN(n6051) );
  NR4D0 U2199 ( .A1(n6054), .A2(n6053), .A3(n6052), .A4(n6051), .ZN(n6076) );
  AOI22D0 U2200 ( .A1(n6933), .A2(\mem[97][6] ), .B1(n6916), .B2(\mem[85][6] ), 
        .ZN(n6058) );
  AOI22D0 U2201 ( .A1(n6935), .A2(\mem[127][6] ), .B1(n6915), .B2(\mem[77][6] ), .ZN(n6057) );
  AOI22D0 U2202 ( .A1(n6979), .A2(\mem[78][6] ), .B1(n6913), .B2(\mem[91][6] ), 
        .ZN(n6056) );
  AOI22D0 U2203 ( .A1(n6969), .A2(\mem[82][6] ), .B1(n6888), .B2(\mem[64][6] ), 
        .ZN(n6055) );
  ND4D0 U2204 ( .A1(n6058), .A2(n6057), .A3(n6056), .A4(n6055), .ZN(n6074) );
  AOI22D0 U2205 ( .A1(n6989), .A2(\mem[70][6] ), .B1(n6296), .B2(\mem[93][6] ), 
        .ZN(n6062) );
  AOI22D0 U2206 ( .A1(n6733), .A2(\mem[122][6] ), .B1(n6680), .B2(\mem[95][6] ), .ZN(n6061) );
  AOI22D0 U2207 ( .A1(n6936), .A2(\mem[81][6] ), .B1(n6982), .B2(\mem[66][6] ), 
        .ZN(n6060) );
  AOI22D0 U2208 ( .A1(n6842), .A2(\mem[90][6] ), .B1(n6847), .B2(\mem[89][6] ), 
        .ZN(n6059) );
  ND4D0 U2209 ( .A1(n6062), .A2(n6061), .A3(n6060), .A4(n6059), .ZN(n6073) );
  AOI22D0 U2210 ( .A1(n6325), .A2(\mem[75][6] ), .B1(n6993), .B2(\mem[117][6] ), .ZN(n6066) );
  AOI22D0 U2211 ( .A1(n6892), .A2(\mem[108][6] ), .B1(n6902), .B2(
        \mem[101][6] ), .ZN(n6065) );
  AOI22D0 U2212 ( .A1(n6970), .A2(\mem[80][6] ), .B1(n6923), .B2(\mem[98][6] ), 
        .ZN(n6063) );
  ND4D0 U2213 ( .A1(n6066), .A2(n6065), .A3(n6064), .A4(n6063), .ZN(n6072) );
  AOI22D0 U2214 ( .A1(n6165), .A2(\mem[110][6] ), .B1(n6990), .B2(\mem[76][6] ), .ZN(n6070) );
  AOI22D0 U2215 ( .A1(n6658), .A2(\mem[114][6] ), .B1(n6869), .B2(
        \mem[113][6] ), .ZN(n6069) );
  AOI22D0 U2216 ( .A1(n6829), .A2(\mem[102][6] ), .B1(n6957), .B2(
        \mem[121][6] ), .ZN(n6068) );
  AOI22D0 U2217 ( .A1(n6981), .A2(\mem[124][6] ), .B1(n6814), .B2(\mem[65][6] ), .ZN(n6067) );
  ND4D0 U2218 ( .A1(n6070), .A2(n6069), .A3(n6068), .A4(n6067), .ZN(n6071) );
  NR4D0 U2219 ( .A1(n6074), .A2(n6073), .A3(n6072), .A4(n6071), .ZN(n6075) );
  CKND2D0 U2220 ( .A1(n6076), .A2(n6075), .ZN(n6163) );
  AOI22D0 U2221 ( .A1(n6928), .A2(\mem[7][6] ), .B1(n6680), .B2(\mem[31][6] ), 
        .ZN(n6080) );
  AOI22D0 U2222 ( .A1(n6658), .A2(\mem[50][6] ), .B1(n6563), .B2(\mem[8][6] ), 
        .ZN(n6079) );
  AOI22D0 U2223 ( .A1(n6860), .A2(\mem[35][6] ), .B1(n6988), .B2(\mem[63][6] ), 
        .ZN(n6078) );
  AOI22D0 U2224 ( .A1(n6614), .A2(\mem[22][6] ), .B1(n6964), .B2(\mem[30][6] ), 
        .ZN(n6077) );
  AOI22D0 U2225 ( .A1(n6989), .A2(\mem[6][6] ), .B1(n6882), .B2(\mem[15][6] ), 
        .ZN(n6084) );
  AOI22D0 U2226 ( .A1(n6905), .A2(\mem[59][6] ), .B1(n6933), .B2(\mem[33][6] ), 
        .ZN(n6083) );
  AOI22D0 U2227 ( .A1(n6179), .A2(\mem[47][6] ), .B1(n6874), .B2(\mem[42][6] ), 
        .ZN(n6082) );
  AOI22D0 U2228 ( .A1(n6936), .A2(\mem[17][6] ), .B1(n6789), .B2(\mem[62][6] ), 
        .ZN(n6081) );
  ND4D0 U2229 ( .A1(n6084), .A2(n6083), .A3(n6082), .A4(n6081), .ZN(n6095) );
  AOI22D0 U2230 ( .A1(n6165), .A2(\mem[46][6] ), .B1(n6915), .B2(\mem[13][6] ), 
        .ZN(n6088) );
  AOI22D0 U2231 ( .A1(n6859), .A2(\mem[52][6] ), .B1(n6804), .B2(\mem[19][6] ), 
        .ZN(n6086) );
  AOI22D0 U2232 ( .A1(n6870), .A2(\mem[60][6] ), .B1(n6749), .B2(\mem[43][6] ), 
        .ZN(n6085) );
  ND4D0 U2233 ( .A1(n6088), .A2(n6087), .A3(n6086), .A4(n6085), .ZN(n6094) );
  AOI22D0 U2234 ( .A1(n6934), .A2(\mem[24][6] ), .B1(n6912), .B2(\mem[56][6] ), 
        .ZN(n6092) );
  AOI22D0 U2235 ( .A1(n6892), .A2(\mem[44][6] ), .B1(n6926), .B2(\mem[1][6] ), 
        .ZN(n6091) );
  AOI22D0 U2236 ( .A1(n6925), .A2(\mem[45][6] ), .B1(n6174), .B2(\mem[54][6] ), 
        .ZN(n6090) );
  AOI22D0 U2237 ( .A1(n6889), .A2(\mem[28][6] ), .B1(n6639), .B2(\mem[39][6] ), 
        .ZN(n6089) );
  ND4D0 U2238 ( .A1(n6092), .A2(n6091), .A3(n6090), .A4(n6089), .ZN(n6093) );
  NR4D0 U2239 ( .A1(n6096), .A2(n6095), .A3(n6094), .A4(n6093), .ZN(n6118) );
  AOI22D0 U2240 ( .A1(n6325), .A2(\mem[11][6] ), .B1(n6993), .B2(\mem[53][6] ), 
        .ZN(n6100) );
  AOI22D0 U2241 ( .A1(n6971), .A2(\mem[38][6] ), .B1(n6774), .B2(\mem[49][6] ), 
        .ZN(n6099) );
  AOI22D0 U2242 ( .A1(n6863), .A2(\mem[55][6] ), .B1(n6955), .B2(\mem[21][6] ), 
        .ZN(n6098) );
  AOI22D0 U2243 ( .A1(n6901), .A2(\mem[9][6] ), .B1(n6924), .B2(\mem[32][6] ), 
        .ZN(n6097) );
  ND4D0 U2244 ( .A1(n6100), .A2(n6099), .A3(n6098), .A4(n6097), .ZN(n6116) );
  AOI22D0 U2245 ( .A1(n6902), .A2(\mem[37][6] ), .B1(n6990), .B2(\mem[12][6] ), 
        .ZN(n6104) );
  AOI22D0 U2246 ( .A1(n6835), .A2(\mem[4][6] ), .B1(n6923), .B2(\mem[34][6] ), 
        .ZN(n6103) );
  AOI22D0 U2247 ( .A1(n6891), .A2(\mem[26][6] ), .B1(n6913), .B2(\mem[27][6] ), 
        .ZN(n6102) );
  AOI22D0 U2248 ( .A1(n6991), .A2(\mem[20][6] ), .B1(n6698), .B2(\mem[2][6] ), 
        .ZN(n6101) );
  ND4D0 U2249 ( .A1(n6104), .A2(n6103), .A3(n6102), .A4(n6101), .ZN(n6115) );
  AOI22D0 U2250 ( .A1(n6759), .A2(\mem[14][6] ), .B1(n6491), .B2(\mem[51][6] ), 
        .ZN(n6107) );
  AOI22D0 U2251 ( .A1(n6773), .A2(\mem[36][6] ), .B1(n6954), .B2(\mem[10][6] ), 
        .ZN(n6106) );
  AOI22D0 U2252 ( .A1(n6542), .A2(\mem[18][6] ), .B1(n6754), .B2(\mem[5][6] ), 
        .ZN(n6105) );
  ND4D0 U2253 ( .A1(n6108), .A2(n6107), .A3(n6106), .A4(n6105), .ZN(n6114) );
  AOI22D0 U2254 ( .A1(n6883), .A2(\mem[48][6] ), .B1(n6847), .B2(\mem[25][6] ), 
        .ZN(n6112) );
  AOI22D0 U2255 ( .A1(n6881), .A2(\mem[16][6] ), .B1(n6879), .B2(\mem[58][6] ), 
        .ZN(n6111) );
  AOI22D0 U2256 ( .A1(n6980), .A2(\mem[61][6] ), .B1(n6957), .B2(\mem[57][6] ), 
        .ZN(n6110) );
  AOI22D0 U2257 ( .A1(n6888), .A2(\mem[0][6] ), .B1(n6995), .B2(\mem[23][6] ), 
        .ZN(n6109) );
  ND4D0 U2258 ( .A1(n6112), .A2(n6111), .A3(n6110), .A4(n6109), .ZN(n6113) );
  NR4D0 U2259 ( .A1(n6116), .A2(n6115), .A3(n6114), .A4(n6113), .ZN(n6117) );
  AOI22D0 U2260 ( .A1(n6728), .A2(\mem[244][6] ), .B1(n6174), .B2(
        \mem[246][6] ), .ZN(n6122) );
  AOI22D0 U2261 ( .A1(n6179), .A2(\mem[239][6] ), .B1(n6542), .B2(
        \mem[210][6] ), .ZN(n6121) );
  AOI22D0 U2262 ( .A1(n6970), .A2(\mem[208][6] ), .B1(n6748), .B2(
        \mem[233][6] ), .ZN(n6120) );
  AOI22D0 U2263 ( .A1(n6980), .A2(\mem[253][6] ), .B1(n6989), .B2(
        \mem[198][6] ), .ZN(n6119) );
  ND4D0 U2264 ( .A1(n6122), .A2(n6121), .A3(n6120), .A4(n6119), .ZN(n6138) );
  AOI22D0 U2265 ( .A1(n6883), .A2(\mem[240][6] ), .B1(n6707), .B2(
        \mem[215][6] ), .ZN(n6126) );
  AOI22D0 U2266 ( .A1(n6994), .A2(\mem[254][6] ), .B1(n6563), .B2(
        \mem[200][6] ), .ZN(n6125) );
  AOI22D0 U2267 ( .A1(n6889), .A2(\mem[220][6] ), .B1(n6990), .B2(
        \mem[204][6] ), .ZN(n6124) );
  ND4D0 U2268 ( .A1(n6126), .A2(n6125), .A3(n6124), .A4(n6123), .ZN(n6137) );
  AOI22D0 U2269 ( .A1(n6928), .A2(\mem[199][6] ), .B1(n6924), .B2(
        \mem[224][6] ), .ZN(n6130) );
  AOI22D0 U2270 ( .A1(n6955), .A2(\mem[213][6] ), .B1(n6957), .B2(
        \mem[249][6] ), .ZN(n6129) );
  AOI22D0 U2271 ( .A1(n6934), .A2(\mem[216][6] ), .B1(n6913), .B2(
        \mem[219][6] ), .ZN(n6128) );
  AOI22D0 U2272 ( .A1(n6981), .A2(\mem[252][6] ), .B1(n6912), .B2(
        \mem[248][6] ), .ZN(n6127) );
  ND4D0 U2273 ( .A1(n6130), .A2(n6129), .A3(n6128), .A4(n6127), .ZN(n6136) );
  AOI22D0 U2274 ( .A1(n6959), .A2(\mem[195][6] ), .B1(n6933), .B2(
        \mem[225][6] ), .ZN(n6134) );
  AOI22D0 U2275 ( .A1(n6165), .A2(\mem[238][6] ), .B1(n6829), .B2(
        \mem[230][6] ), .ZN(n6133) );
  AOI22D0 U2276 ( .A1(n6979), .A2(\mem[206][6] ), .B1(n6902), .B2(
        \mem[229][6] ), .ZN(n6132) );
  AOI22D0 U2277 ( .A1(n6760), .A2(\mem[237][6] ), .B1(n6882), .B2(
        \mem[207][6] ), .ZN(n6131) );
  ND4D0 U2278 ( .A1(n6134), .A2(n6133), .A3(n6132), .A4(n6131), .ZN(n6135) );
  NR4D0 U2279 ( .A1(n6138), .A2(n6137), .A3(n6136), .A4(n6135), .ZN(n6160) );
  AOI22D0 U2280 ( .A1(n6976), .A2(\mem[226][6] ), .B1(n6956), .B2(
        \mem[232][6] ), .ZN(n6142) );
  AOI22D0 U2281 ( .A1(n6680), .A2(\mem[223][6] ), .B1(n6993), .B2(
        \mem[245][6] ), .ZN(n6141) );
  AOI22D0 U2282 ( .A1(n6809), .A2(\mem[201][6] ), .B1(n6936), .B2(
        \mem[209][6] ), .ZN(n6140) );
  AOI22D0 U2283 ( .A1(n6614), .A2(\mem[214][6] ), .B1(n6888), .B2(
        \mem[192][6] ), .ZN(n6139) );
  ND4D0 U2284 ( .A1(n6142), .A2(n6141), .A3(n6140), .A4(n6139), .ZN(n6158) );
  AOI22D0 U2285 ( .A1(n6747), .A2(\mem[212][6] ), .B1(n6879), .B2(
        \mem[250][6] ), .ZN(n6146) );
  AOI22D0 U2286 ( .A1(n6890), .A2(\mem[228][6] ), .B1(n6835), .B2(
        \mem[196][6] ), .ZN(n6145) );
  AOI22D0 U2287 ( .A1(n6749), .A2(\mem[235][6] ), .B1(n6880), .B2(
        \mem[203][6] ), .ZN(n6143) );
  ND4D0 U2288 ( .A1(n6146), .A2(n6145), .A3(n6144), .A4(n6143), .ZN(n6157) );
  AOI22D0 U2289 ( .A1(n6860), .A2(\mem[227][6] ), .B1(n6954), .B2(
        \mem[202][6] ), .ZN(n6150) );
  AOI22D0 U2290 ( .A1(n6658), .A2(\mem[242][6] ), .B1(n6982), .B2(
        \mem[194][6] ), .ZN(n6149) );
  AOI22D0 U2291 ( .A1(n6639), .A2(\mem[231][6] ), .B1(n6804), .B2(
        \mem[211][6] ), .ZN(n6148) );
  AOI22D0 U2292 ( .A1(n6892), .A2(\mem[236][6] ), .B1(n6914), .B2(
        \mem[197][6] ), .ZN(n6147) );
  ND4D0 U2293 ( .A1(n6150), .A2(n6149), .A3(n6148), .A4(n6147), .ZN(n6156) );
  AOI22D0 U2294 ( .A1(n6814), .A2(\mem[193][6] ), .B1(n6296), .B2(
        \mem[221][6] ), .ZN(n6154) );
  AOI22D0 U2295 ( .A1(n6891), .A2(\mem[218][6] ), .B1(n6774), .B2(
        \mem[241][6] ), .ZN(n6153) );
  AOI22D0 U2296 ( .A1(n6905), .A2(\mem[251][6] ), .B1(n6964), .B2(
        \mem[222][6] ), .ZN(n6152) );
  AOI22D0 U2297 ( .A1(n6491), .A2(\mem[243][6] ), .B1(n6847), .B2(
        \mem[217][6] ), .ZN(n6151) );
  NR4D0 U2298 ( .A1(n6158), .A2(n6157), .A3(n6156), .A4(n6155), .ZN(n6159) );
  AOI21D0 U2299 ( .A1(n6160), .A2(n6159), .B(n6945), .ZN(n6161) );
  AOI211D0 U2300 ( .A1(n6164), .A2(n6163), .B(n6162), .C(n6161), .ZN(n6190) );
  AOI22D0 U2301 ( .A1(n6165), .A2(\mem[174][6] ), .B1(n6842), .B2(
        \mem[154][6] ), .ZN(n6169) );
  AOI22D0 U2302 ( .A1(n6991), .A2(\mem[148][6] ), .B1(n6983), .B2(
        \mem[176][6] ), .ZN(n6168) );
  AOI22D0 U2303 ( .A1(n6749), .A2(\mem[171][6] ), .B1(n6935), .B2(
        \mem[191][6] ), .ZN(n6167) );
  AOI22D0 U2304 ( .A1(n6969), .A2(\mem[146][6] ), .B1(n6993), .B2(
        \mem[181][6] ), .ZN(n6166) );
  ND4D0 U2305 ( .A1(n6169), .A2(n6168), .A3(n6167), .A4(n6166), .ZN(n6187) );
  AOI22D0 U2306 ( .A1(n6981), .A2(\mem[188][6] ), .B1(n6789), .B2(
        \mem[190][6] ), .ZN(n6173) );
  AOI22D0 U2307 ( .A1(n6933), .A2(\mem[161][6] ), .B1(n6296), .B2(
        \mem[157][6] ), .ZN(n6172) );
  AOI22D0 U2308 ( .A1(n6905), .A2(\mem[187][6] ), .B1(n6901), .B2(
        \mem[137][6] ), .ZN(n6171) );
  AOI22D0 U2309 ( .A1(n6814), .A2(\mem[129][6] ), .B1(n6995), .B2(
        \mem[151][6] ), .ZN(n6170) );
  ND4D0 U2310 ( .A1(n6173), .A2(n6172), .A3(n6171), .A4(n6170), .ZN(n6186) );
  AOI22D0 U2311 ( .A1(n6874), .A2(\mem[170][6] ), .B1(n6680), .B2(
        \mem[159][6] ), .ZN(n6178) );
  AOI22D0 U2312 ( .A1(n6325), .A2(\mem[139][6] ), .B1(n6913), .B2(
        \mem[155][6] ), .ZN(n6177) );
  AOI22D0 U2313 ( .A1(n6803), .A2(\mem[183][6] ), .B1(n6174), .B2(
        \mem[182][6] ), .ZN(n6176) );
  AOI22D0 U2314 ( .A1(n6829), .A2(\mem[166][6] ), .B1(n6698), .B2(
        \mem[130][6] ), .ZN(n6175) );
  ND4D0 U2315 ( .A1(n6178), .A2(n6177), .A3(n6176), .A4(n6175), .ZN(n6185) );
  AOI22D0 U2316 ( .A1(n6802), .A2(\mem[152][6] ), .B1(n6733), .B2(
        \mem[186][6] ), .ZN(n6183) );
  AOI22D0 U2317 ( .A1(n6179), .A2(\mem[175][6] ), .B1(n6639), .B2(
        \mem[167][6] ), .ZN(n6182) );
  AOI22D0 U2318 ( .A1(n6860), .A2(\mem[163][6] ), .B1(n6923), .B2(
        \mem[162][6] ), .ZN(n6180) );
  ND4D0 U2319 ( .A1(n6183), .A2(n6182), .A3(n6181), .A4(n6180), .ZN(n6184) );
  NR4D0 U2320 ( .A1(n6187), .A2(n6186), .A3(n6185), .A4(n6184), .ZN(n6189) );
  AOI32D0 U2321 ( .A1(n6191), .A2(n6190), .A3(n6189), .B1(n6188), .B2(n6190), 
        .ZN(dout[6]) );
  AOI22D0 U2322 ( .A1(n6989), .A2(\mem[70][7] ), .B1(n6991), .B2(\mem[84][7] ), 
        .ZN(n6195) );
  AOI22D0 U2323 ( .A1(n6325), .A2(\mem[75][7] ), .B1(n6862), .B2(\mem[104][7] ), .ZN(n6194) );
  AOI22D0 U2324 ( .A1(n6809), .A2(\mem[73][7] ), .B1(n6837), .B2(\mem[79][7] ), 
        .ZN(n6193) );
  AOI22D0 U2325 ( .A1(n6922), .A2(\mem[93][7] ), .B1(n6993), .B2(\mem[117][7] ), .ZN(n6192) );
  ND4D0 U2326 ( .A1(n6195), .A2(n6194), .A3(n6193), .A4(n6192), .ZN(n6211) );
  AOI22D0 U2327 ( .A1(n6967), .A2(\mem[103][7] ), .B1(n6982), .B2(\mem[66][7] ), .ZN(n6199) );
  AOI22D0 U2328 ( .A1(n6926), .A2(\mem[65][7] ), .B1(n6873), .B2(\mem[94][7] ), 
        .ZN(n6198) );
  AOI22D0 U2329 ( .A1(n6891), .A2(\mem[90][7] ), .B1(n6992), .B2(\mem[118][7] ), .ZN(n6197) );
  AOI22D0 U2330 ( .A1(n6959), .A2(\mem[67][7] ), .B1(n6916), .B2(\mem[85][7] ), 
        .ZN(n6196) );
  ND4D0 U2331 ( .A1(n6199), .A2(n6198), .A3(n6197), .A4(n6196), .ZN(n6210) );
  AOI22D0 U2332 ( .A1(n6860), .A2(\mem[99][7] ), .B1(n6969), .B2(\mem[82][7] ), 
        .ZN(n6202) );
  AOI22D0 U2333 ( .A1(n6890), .A2(\mem[100][7] ), .B1(n6888), .B2(\mem[64][7] ), .ZN(n6201) );
  AOI22D0 U2334 ( .A1(n6953), .A2(\mem[111][7] ), .B1(n6935), .B2(
        \mem[127][7] ), .ZN(n6200) );
  ND4D0 U2335 ( .A1(n6203), .A2(n6202), .A3(n6201), .A4(n6200), .ZN(n6209) );
  AOI22D0 U2336 ( .A1(n6980), .A2(\mem[125][7] ), .B1(n6892), .B2(
        \mem[108][7] ), .ZN(n6207) );
  AOI22D0 U2337 ( .A1(n6927), .A2(\mem[89][7] ), .B1(n6994), .B2(\mem[126][7] ), .ZN(n6206) );
  AOI22D0 U2338 ( .A1(n6928), .A2(\mem[71][7] ), .B1(n6979), .B2(\mem[78][7] ), 
        .ZN(n6205) );
  AOI22D0 U2339 ( .A1(n6952), .A2(\mem[86][7] ), .B1(n6563), .B2(\mem[72][7] ), 
        .ZN(n6204) );
  ND4D0 U2340 ( .A1(n6207), .A2(n6206), .A3(n6205), .A4(n6204), .ZN(n6208) );
  NR4D0 U2341 ( .A1(n6211), .A2(n6210), .A3(n6209), .A4(n6208), .ZN(n6365) );
  AOI22D0 U2342 ( .A1(n6991), .A2(\mem[148][7] ), .B1(n6837), .B2(
        \mem[143][7] ), .ZN(n6215) );
  AOI22D0 U2343 ( .A1(n6773), .A2(\mem[164][7] ), .B1(n6993), .B2(
        \mem[181][7] ), .ZN(n6214) );
  AOI22D0 U2344 ( .A1(n6868), .A2(\mem[171][7] ), .B1(n6871), .B2(
        \mem[185][7] ), .ZN(n6213) );
  AOI22D0 U2345 ( .A1(n6860), .A2(\mem[163][7] ), .B1(n6970), .B2(
        \mem[144][7] ), .ZN(n6212) );
  ND4D0 U2346 ( .A1(n6215), .A2(n6214), .A3(n6213), .A4(n6212), .ZN(n6231) );
  AOI22D0 U2347 ( .A1(n6542), .A2(\mem[146][7] ), .B1(n6891), .B2(
        \mem[154][7] ), .ZN(n6219) );
  AOI22D0 U2348 ( .A1(n6982), .A2(\mem[130][7] ), .B1(n6992), .B2(
        \mem[182][7] ), .ZN(n6217) );
  AOI22D0 U2349 ( .A1(n6760), .A2(\mem[173][7] ), .B1(n6563), .B2(
        \mem[136][7] ), .ZN(n6216) );
  ND4D0 U2350 ( .A1(n6219), .A2(n6218), .A3(n6217), .A4(n6216), .ZN(n6230) );
  AOI22D0 U2351 ( .A1(n6889), .A2(\mem[156][7] ), .B1(n6873), .B2(
        \mem[158][7] ), .ZN(n6223) );
  AOI22D0 U2352 ( .A1(n6859), .A2(\mem[180][7] ), .B1(n6935), .B2(
        \mem[191][7] ), .ZN(n6222) );
  AOI22D0 U2353 ( .A1(n6983), .A2(\mem[176][7] ), .B1(n6804), .B2(
        \mem[147][7] ), .ZN(n6221) );
  AOI22D0 U2354 ( .A1(n6981), .A2(\mem[188][7] ), .B1(n6979), .B2(
        \mem[142][7] ), .ZN(n6220) );
  ND4D0 U2355 ( .A1(n6223), .A2(n6222), .A3(n6221), .A4(n6220), .ZN(n6229) );
  AOI22D0 U2356 ( .A1(n6879), .A2(\mem[186][7] ), .B1(n6966), .B2(
        \mem[178][7] ), .ZN(n6227) );
  AOI22D0 U2357 ( .A1(n6847), .A2(\mem[153][7] ), .B1(n6955), .B2(
        \mem[149][7] ), .ZN(n6226) );
  AOI22D0 U2358 ( .A1(n6959), .A2(\mem[131][7] ), .B1(n6995), .B2(
        \mem[151][7] ), .ZN(n6225) );
  AOI22D0 U2359 ( .A1(n6680), .A2(\mem[159][7] ), .B1(n6994), .B2(
        \mem[190][7] ), .ZN(n6224) );
  ND4D0 U2360 ( .A1(n6227), .A2(n6226), .A3(n6225), .A4(n6224), .ZN(n6228) );
  NR4D0 U2361 ( .A1(n6231), .A2(n6230), .A3(n6229), .A4(n6228), .ZN(n6253) );
  AOI22D0 U2362 ( .A1(n6917), .A2(\mem[174][7] ), .B1(n6980), .B2(
        \mem[189][7] ), .ZN(n6235) );
  AOI22D0 U2363 ( .A1(n6905), .A2(\mem[187][7] ), .B1(n6861), .B2(
        \mem[132][7] ), .ZN(n6234) );
  AOI22D0 U2364 ( .A1(n6967), .A2(\mem[167][7] ), .B1(n6912), .B2(
        \mem[184][7] ), .ZN(n6233) );
  AOI22D0 U2365 ( .A1(n6888), .A2(\mem[128][7] ), .B1(n6990), .B2(
        \mem[140][7] ), .ZN(n6232) );
  ND4D0 U2366 ( .A1(n6235), .A2(n6234), .A3(n6233), .A4(n6232), .ZN(n6251) );
  AOI22D0 U2367 ( .A1(n6977), .A2(\mem[161][7] ), .B1(n6923), .B2(
        \mem[162][7] ), .ZN(n6238) );
  AOI22D0 U2368 ( .A1(n6892), .A2(\mem[172][7] ), .B1(n6915), .B2(
        \mem[141][7] ), .ZN(n6237) );
  AOI22D0 U2369 ( .A1(n6325), .A2(\mem[139][7] ), .B1(n6958), .B2(
        \mem[145][7] ), .ZN(n6236) );
  ND4D0 U2370 ( .A1(n6239), .A2(n6238), .A3(n6237), .A4(n6236), .ZN(n6250) );
  AOI22D0 U2371 ( .A1(n6614), .A2(\mem[150][7] ), .B1(n6989), .B2(
        \mem[134][7] ), .ZN(n6243) );
  AOI22D0 U2372 ( .A1(n6926), .A2(\mem[129][7] ), .B1(n6956), .B2(
        \mem[168][7] ), .ZN(n6242) );
  AOI22D0 U2373 ( .A1(n6953), .A2(\mem[175][7] ), .B1(n6902), .B2(
        \mem[165][7] ), .ZN(n6241) );
  AOI22D0 U2374 ( .A1(n6790), .A2(\mem[155][7] ), .B1(n6903), .B2(
        \mem[179][7] ), .ZN(n6240) );
  ND4D0 U2375 ( .A1(n6243), .A2(n6242), .A3(n6241), .A4(n6240), .ZN(n6249) );
  AOI22D0 U2376 ( .A1(n6914), .A2(\mem[133][7] ), .B1(n6924), .B2(
        \mem[160][7] ), .ZN(n6247) );
  AOI22D0 U2377 ( .A1(n6971), .A2(\mem[166][7] ), .B1(n6954), .B2(
        \mem[138][7] ), .ZN(n6246) );
  AOI22D0 U2378 ( .A1(n6874), .A2(\mem[170][7] ), .B1(n6296), .B2(
        \mem[157][7] ), .ZN(n6245) );
  AOI22D0 U2379 ( .A1(n6934), .A2(\mem[152][7] ), .B1(n6809), .B2(
        \mem[137][7] ), .ZN(n6244) );
  ND4D0 U2380 ( .A1(n6247), .A2(n6246), .A3(n6245), .A4(n6244), .ZN(n6248) );
  NR4D0 U2381 ( .A1(n6251), .A2(n6250), .A3(n6249), .A4(n6248), .ZN(n6252) );
  CKND2D0 U2382 ( .A1(n6253), .A2(n6252), .ZN(n6342) );
  AOI22D0 U2383 ( .A1(n6861), .A2(\mem[4][7] ), .B1(n6874), .B2(\mem[42][7] ), 
        .ZN(n6257) );
  AOI22D0 U2384 ( .A1(n6981), .A2(\mem[60][7] ), .B1(n6873), .B2(\mem[30][7] ), 
        .ZN(n6256) );
  AOI22D0 U2385 ( .A1(n6658), .A2(\mem[50][7] ), .B1(n6990), .B2(\mem[12][7] ), 
        .ZN(n6255) );
  ND4D0 U2386 ( .A1(n6257), .A2(n6256), .A3(n6255), .A4(n6254), .ZN(n6273) );
  AOI22D0 U2387 ( .A1(n6836), .A2(\mem[10][7] ), .B1(n6563), .B2(\mem[8][7] ), 
        .ZN(n6261) );
  AOI22D0 U2388 ( .A1(n6890), .A2(\mem[36][7] ), .B1(n6979), .B2(\mem[14][7] ), 
        .ZN(n6260) );
  AOI22D0 U2389 ( .A1(n6989), .A2(\mem[6][7] ), .B1(n6958), .B2(\mem[17][7] ), 
        .ZN(n6259) );
  AOI22D0 U2390 ( .A1(n6659), .A2(\mem[53][7] ), .B1(n6915), .B2(\mem[13][7] ), 
        .ZN(n6258) );
  ND4D0 U2391 ( .A1(n6261), .A2(n6260), .A3(n6259), .A4(n6258), .ZN(n6272) );
  AOI22D0 U2392 ( .A1(n6969), .A2(\mem[18][7] ), .B1(n6847), .B2(\mem[25][7] ), 
        .ZN(n6265) );
  AOI22D0 U2393 ( .A1(n6829), .A2(\mem[38][7] ), .B1(n6968), .B2(\mem[41][7] ), 
        .ZN(n6264) );
  AOI22D0 U2394 ( .A1(n6953), .A2(\mem[47][7] ), .B1(n6680), .B2(\mem[31][7] ), 
        .ZN(n6263) );
  AOI22D0 U2395 ( .A1(n6934), .A2(\mem[24][7] ), .B1(n6956), .B2(\mem[40][7] ), 
        .ZN(n6262) );
  ND4D0 U2396 ( .A1(n6265), .A2(n6264), .A3(n6263), .A4(n6262), .ZN(n6271) );
  AOI22D0 U2397 ( .A1(n6892), .A2(\mem[44][7] ), .B1(n6935), .B2(\mem[63][7] ), 
        .ZN(n6269) );
  AOI22D0 U2398 ( .A1(n6491), .A2(\mem[51][7] ), .B1(n6995), .B2(\mem[23][7] ), 
        .ZN(n6268) );
  AOI22D0 U2399 ( .A1(n6891), .A2(\mem[26][7] ), .B1(n6913), .B2(\mem[27][7] ), 
        .ZN(n6267) );
  AOI22D0 U2400 ( .A1(n6863), .A2(\mem[55][7] ), .B1(n6957), .B2(\mem[57][7] ), 
        .ZN(n6266) );
  ND4D0 U2401 ( .A1(n6269), .A2(n6268), .A3(n6267), .A4(n6266), .ZN(n6270) );
  NR4D0 U2402 ( .A1(n6273), .A2(n6272), .A3(n6271), .A4(n6270), .ZN(n6295) );
  AOI22D0 U2403 ( .A1(n6914), .A2(\mem[5][7] ), .B1(n6901), .B2(\mem[9][7] ), 
        .ZN(n6277) );
  AOI22D0 U2404 ( .A1(n6959), .A2(\mem[3][7] ), .B1(n6902), .B2(\mem[37][7] ), 
        .ZN(n6276) );
  AOI22D0 U2405 ( .A1(n6904), .A2(\mem[19][7] ), .B1(n6869), .B2(\mem[49][7] ), 
        .ZN(n6274) );
  ND4D0 U2406 ( .A1(n6277), .A2(n6276), .A3(n6275), .A4(n6274), .ZN(n6293) );
  AOI22D0 U2407 ( .A1(n6905), .A2(\mem[59][7] ), .B1(n6991), .B2(\mem[20][7] ), 
        .ZN(n6281) );
  AOI22D0 U2408 ( .A1(n6860), .A2(\mem[35][7] ), .B1(n6881), .B2(\mem[16][7] ), 
        .ZN(n6280) );
  AOI22D0 U2409 ( .A1(n6325), .A2(\mem[11][7] ), .B1(n6296), .B2(\mem[29][7] ), 
        .ZN(n6279) );
  AOI22D0 U2410 ( .A1(n6917), .A2(\mem[46][7] ), .B1(n6928), .B2(\mem[7][7] ), 
        .ZN(n6278) );
  ND4D0 U2411 ( .A1(n6281), .A2(n6280), .A3(n6279), .A4(n6278), .ZN(n6292) );
  AOI22D0 U2412 ( .A1(n6888), .A2(\mem[0][7] ), .B1(n6924), .B2(\mem[32][7] ), 
        .ZN(n6285) );
  AOI22D0 U2413 ( .A1(n6925), .A2(\mem[45][7] ), .B1(n6992), .B2(\mem[54][7] ), 
        .ZN(n6284) );
  AOI22D0 U2414 ( .A1(n6976), .A2(\mem[34][7] ), .B1(n6728), .B2(\mem[52][7] ), 
        .ZN(n6283) );
  AOI22D0 U2415 ( .A1(n6980), .A2(\mem[61][7] ), .B1(n6994), .B2(\mem[62][7] ), 
        .ZN(n6282) );
  AOI22D0 U2416 ( .A1(n6784), .A2(\mem[28][7] ), .B1(n6983), .B2(\mem[48][7] ), 
        .ZN(n6289) );
  AOI22D0 U2417 ( .A1(n6933), .A2(\mem[33][7] ), .B1(n6837), .B2(\mem[15][7] ), 
        .ZN(n6288) );
  AOI22D0 U2418 ( .A1(n6749), .A2(\mem[43][7] ), .B1(n6952), .B2(\mem[22][7] ), 
        .ZN(n6287) );
  AOI22D0 U2419 ( .A1(n6814), .A2(\mem[1][7] ), .B1(n6912), .B2(\mem[56][7] ), 
        .ZN(n6286) );
  ND4D0 U2420 ( .A1(n6289), .A2(n6288), .A3(n6287), .A4(n6286), .ZN(n6290) );
  NR4D0 U2421 ( .A1(n6293), .A2(n6292), .A3(n6291), .A4(n6290), .ZN(n6294) );
  AOI22D0 U2422 ( .A1(n6863), .A2(\mem[247][7] ), .B1(n6658), .B2(
        \mem[242][7] ), .ZN(n6300) );
  AOI22D0 U2423 ( .A1(n6749), .A2(\mem[235][7] ), .B1(n6296), .B2(
        \mem[221][7] ), .ZN(n6298) );
  AOI22D0 U2424 ( .A1(n6959), .A2(\mem[195][7] ), .B1(n6491), .B2(
        \mem[243][7] ), .ZN(n6297) );
  ND4D0 U2425 ( .A1(n6300), .A2(n6299), .A3(n6298), .A4(n6297), .ZN(n6316) );
  AOI22D0 U2426 ( .A1(n6883), .A2(\mem[240][7] ), .B1(n6754), .B2(
        \mem[197][7] ), .ZN(n6304) );
  AOI22D0 U2427 ( .A1(n6926), .A2(\mem[193][7] ), .B1(n6933), .B2(
        \mem[225][7] ), .ZN(n6303) );
  AOI22D0 U2428 ( .A1(n6888), .A2(\mem[192][7] ), .B1(n6901), .B2(
        \mem[201][7] ), .ZN(n6302) );
  AOI22D0 U2429 ( .A1(n6791), .A2(\mem[224][7] ), .B1(n6994), .B2(
        \mem[254][7] ), .ZN(n6301) );
  ND4D0 U2430 ( .A1(n6304), .A2(n6303), .A3(n6302), .A4(n6301), .ZN(n6315) );
  AOI22D0 U2431 ( .A1(n6892), .A2(\mem[236][7] ), .B1(n6733), .B2(
        \mem[250][7] ), .ZN(n6308) );
  AOI22D0 U2432 ( .A1(n6980), .A2(\mem[253][7] ), .B1(n6871), .B2(
        \mem[249][7] ), .ZN(n6307) );
  AOI22D0 U2433 ( .A1(n6991), .A2(\mem[212][7] ), .B1(n6837), .B2(
        \mem[207][7] ), .ZN(n6306) );
  AOI22D0 U2434 ( .A1(n6927), .A2(\mem[217][7] ), .B1(n6958), .B2(
        \mem[209][7] ), .ZN(n6305) );
  ND4D0 U2435 ( .A1(n6308), .A2(n6307), .A3(n6306), .A4(n6305), .ZN(n6314) );
  AOI22D0 U2436 ( .A1(n6928), .A2(\mem[199][7] ), .B1(n6891), .B2(
        \mem[218][7] ), .ZN(n6312) );
  AOI22D0 U2437 ( .A1(n6971), .A2(\mem[230][7] ), .B1(n6935), .B2(
        \mem[255][7] ), .ZN(n6311) );
  AOI22D0 U2438 ( .A1(n6953), .A2(\mem[239][7] ), .B1(n6912), .B2(
        \mem[248][7] ), .ZN(n6310) );
  AOI22D0 U2439 ( .A1(n6916), .A2(\mem[213][7] ), .B1(n6954), .B2(
        \mem[202][7] ), .ZN(n6309) );
  ND4D0 U2440 ( .A1(n6312), .A2(n6311), .A3(n6310), .A4(n6309), .ZN(n6313) );
  NR4D0 U2441 ( .A1(n6316), .A2(n6315), .A3(n6314), .A4(n6313), .ZN(n6339) );
  AOI22D0 U2442 ( .A1(n6760), .A2(\mem[237][7] ), .B1(n6738), .B2(
        \mem[229][7] ), .ZN(n6319) );
  AOI22D0 U2443 ( .A1(n6968), .A2(\mem[233][7] ), .B1(n6873), .B2(
        \mem[222][7] ), .ZN(n6318) );
  AOI22D0 U2444 ( .A1(n6614), .A2(\mem[214][7] ), .B1(n6728), .B2(
        \mem[244][7] ), .ZN(n6317) );
  ND4D0 U2445 ( .A1(n6320), .A2(n6319), .A3(n6318), .A4(n6317), .ZN(n6337) );
  AOI22D0 U2446 ( .A1(n6905), .A2(\mem[251][7] ), .B1(n6993), .B2(
        \mem[245][7] ), .ZN(n6324) );
  AOI22D0 U2447 ( .A1(n6860), .A2(\mem[227][7] ), .B1(n6906), .B2(
        \mem[204][7] ), .ZN(n6323) );
  AOI22D0 U2448 ( .A1(n6978), .A2(\mem[200][7] ), .B1(n6992), .B2(
        \mem[246][7] ), .ZN(n6322) );
  AOI22D0 U2449 ( .A1(n6870), .A2(\mem[252][7] ), .B1(n6639), .B2(
        \mem[231][7] ), .ZN(n6321) );
  ND4D0 U2450 ( .A1(n6324), .A2(n6323), .A3(n6322), .A4(n6321), .ZN(n6336) );
  AOI22D0 U2451 ( .A1(n6934), .A2(\mem[216][7] ), .B1(n6862), .B2(
        \mem[232][7] ), .ZN(n6329) );
  AOI22D0 U2452 ( .A1(n6976), .A2(\mem[226][7] ), .B1(n6869), .B2(
        \mem[241][7] ), .ZN(n6328) );
  AOI22D0 U2453 ( .A1(n6325), .A2(\mem[203][7] ), .B1(n6861), .B2(
        \mem[196][7] ), .ZN(n6327) );
  AOI22D0 U2454 ( .A1(n6989), .A2(\mem[198][7] ), .B1(n6913), .B2(
        \mem[219][7] ), .ZN(n6326) );
  ND4D0 U2455 ( .A1(n6329), .A2(n6328), .A3(n6327), .A4(n6326), .ZN(n6335) );
  AOI22D0 U2456 ( .A1(n6542), .A2(\mem[210][7] ), .B1(n6874), .B2(
        \mem[234][7] ), .ZN(n6333) );
  AOI22D0 U2457 ( .A1(n6680), .A2(\mem[223][7] ), .B1(n6982), .B2(
        \mem[194][7] ), .ZN(n6332) );
  AOI22D0 U2458 ( .A1(n6917), .A2(\mem[238][7] ), .B1(n6881), .B2(
        \mem[208][7] ), .ZN(n6331) );
  ND4D0 U2459 ( .A1(n6333), .A2(n6332), .A3(n6331), .A4(n6330), .ZN(n6334) );
  NR4D0 U2460 ( .A1(n6337), .A2(n6336), .A3(n6335), .A4(n6334), .ZN(n6338) );
  AOI21D0 U2461 ( .A1(n6339), .A2(n6338), .B(n6945), .ZN(n6340) );
  AOI211D0 U2462 ( .A1(n6951), .A2(n6342), .B(n6341), .C(n6340), .ZN(n6364) );
  AOI22D0 U2463 ( .A1(n6933), .A2(\mem[97][7] ), .B1(n6874), .B2(\mem[106][7] ), .ZN(n6346) );
  AOI22D0 U2464 ( .A1(n6981), .A2(\mem[124][7] ), .B1(n6957), .B2(
        \mem[121][7] ), .ZN(n6344) );
  AOI22D0 U2465 ( .A1(n6917), .A2(\mem[110][7] ), .B1(n6990), .B2(\mem[76][7] ), .ZN(n6343) );
  ND4D0 U2466 ( .A1(n6346), .A2(n6345), .A3(n6344), .A4(n6343), .ZN(n6362) );
  AOI22D0 U2467 ( .A1(n6784), .A2(\mem[92][7] ), .B1(n6903), .B2(\mem[115][7] ), .ZN(n6350) );
  AOI22D0 U2468 ( .A1(n6680), .A2(\mem[95][7] ), .B1(n6995), .B2(\mem[87][7] ), 
        .ZN(n6349) );
  AOI22D0 U2469 ( .A1(n6983), .A2(\mem[112][7] ), .B1(n6923), .B2(\mem[98][7] ), .ZN(n6348) );
  AOI22D0 U2470 ( .A1(n6802), .A2(\mem[88][7] ), .B1(n6829), .B2(\mem[102][7] ), .ZN(n6347) );
  ND4D0 U2471 ( .A1(n6350), .A2(n6349), .A3(n6348), .A4(n6347), .ZN(n6361) );
  AOI22D0 U2472 ( .A1(n6804), .A2(\mem[83][7] ), .B1(n6828), .B2(\mem[120][7] ), .ZN(n6354) );
  AOI22D0 U2473 ( .A1(n6835), .A2(\mem[68][7] ), .B1(n6738), .B2(\mem[101][7] ), .ZN(n6353) );
  AOI22D0 U2474 ( .A1(n6970), .A2(\mem[80][7] ), .B1(n6924), .B2(\mem[96][7] ), 
        .ZN(n6352) );
  AOI22D0 U2475 ( .A1(n6790), .A2(\mem[91][7] ), .B1(n6658), .B2(\mem[114][7] ), .ZN(n6351) );
  ND4D0 U2476 ( .A1(n6354), .A2(n6353), .A3(n6352), .A4(n6351), .ZN(n6360) );
  AOI22D0 U2477 ( .A1(n6836), .A2(\mem[74][7] ), .B1(n6915), .B2(\mem[77][7] ), 
        .ZN(n6358) );
  AOI22D0 U2478 ( .A1(n6879), .A2(\mem[122][7] ), .B1(n6774), .B2(
        \mem[113][7] ), .ZN(n6357) );
  AOI22D0 U2479 ( .A1(n6863), .A2(\mem[119][7] ), .B1(n6936), .B2(\mem[81][7] ), .ZN(n6356) );
  AOI22D0 U2480 ( .A1(n6905), .A2(\mem[123][7] ), .B1(n6728), .B2(
        \mem[116][7] ), .ZN(n6355) );
  ND4D0 U2481 ( .A1(n6358), .A2(n6357), .A3(n6356), .A4(n6355), .ZN(n6359) );
  NR4D0 U2482 ( .A1(n6362), .A2(n6361), .A3(n6360), .A4(n6359), .ZN(n6363) );
  AOI32D0 U2483 ( .A1(n6365), .A2(n6364), .A3(n6363), .B1(n7004), .B2(n6364), 
        .ZN(dout[7]) );
  AOI22D0 U2484 ( .A1(n6959), .A2(\mem[3][2] ), .B1(n6892), .B2(\mem[44][2] ), 
        .ZN(n6368) );
  AOI22D0 U2485 ( .A1(n6889), .A2(\mem[28][2] ), .B1(n6707), .B2(\mem[23][2] ), 
        .ZN(n6367) );
  AOI22D0 U2486 ( .A1(n6861), .A2(\mem[4][2] ), .B1(n6891), .B2(\mem[26][2] ), 
        .ZN(n6366) );
  ND4D0 U2487 ( .A1(n6369), .A2(n6368), .A3(n6367), .A4(n6366), .ZN(n6385) );
  AOI22D0 U2488 ( .A1(n6880), .A2(\mem[11][2] ), .B1(n6760), .B2(\mem[45][2] ), 
        .ZN(n6373) );
  AOI22D0 U2489 ( .A1(n6923), .A2(\mem[34][2] ), .B1(n6804), .B2(\mem[19][2] ), 
        .ZN(n6372) );
  AOI22D0 U2490 ( .A1(n6981), .A2(\mem[60][2] ), .B1(n6733), .B2(\mem[58][2] ), 
        .ZN(n6371) );
  AOI22D0 U2491 ( .A1(n6809), .A2(\mem[9][2] ), .B1(n6935), .B2(\mem[63][2] ), 
        .ZN(n6370) );
  ND4D0 U2492 ( .A1(n6373), .A2(n6372), .A3(n6371), .A4(n6370), .ZN(n6384) );
  AOI22D0 U2493 ( .A1(n6922), .A2(\mem[29][2] ), .B1(n6992), .B2(\mem[54][2] ), 
        .ZN(n6377) );
  AOI22D0 U2494 ( .A1(n6955), .A2(\mem[21][2] ), .B1(n6906), .B2(\mem[12][2] ), 
        .ZN(n6376) );
  AOI22D0 U2495 ( .A1(n6980), .A2(\mem[61][2] ), .B1(n6924), .B2(\mem[32][2] ), 
        .ZN(n6375) );
  AOI22D0 U2496 ( .A1(n6991), .A2(\mem[20][2] ), .B1(n6964), .B2(\mem[30][2] ), 
        .ZN(n6374) );
  ND4D0 U2497 ( .A1(n6377), .A2(n6376), .A3(n6375), .A4(n6374), .ZN(n6383) );
  AOI22D0 U2498 ( .A1(n6883), .A2(\mem[48][2] ), .B1(n6738), .B2(\mem[37][2] ), 
        .ZN(n6381) );
  AOI22D0 U2499 ( .A1(n6979), .A2(\mem[14][2] ), .B1(n5966), .B2(\mem[31][2] ), 
        .ZN(n6380) );
  AOI22D0 U2500 ( .A1(n6874), .A2(\mem[42][2] ), .B1(n6927), .B2(\mem[25][2] ), 
        .ZN(n6379) );
  ND4D0 U2501 ( .A1(n6381), .A2(n6380), .A3(n6379), .A4(n6378), .ZN(n6382) );
  NR4D0 U2502 ( .A1(n6385), .A2(n6384), .A3(n6383), .A4(n6382), .ZN(n6541) );
  AOI22D0 U2503 ( .A1(n6874), .A2(\mem[170][2] ), .B1(n6828), .B2(
        \mem[184][2] ), .ZN(n6389) );
  AOI22D0 U2504 ( .A1(n6983), .A2(\mem[176][2] ), .B1(n6738), .B2(
        \mem[165][2] ), .ZN(n6388) );
  AOI22D0 U2505 ( .A1(n6970), .A2(\mem[144][2] ), .B1(n6837), .B2(
        \mem[143][2] ), .ZN(n6387) );
  AOI22D0 U2506 ( .A1(n6749), .A2(\mem[171][2] ), .B1(n6789), .B2(
        \mem[190][2] ), .ZN(n6386) );
  ND4D0 U2507 ( .A1(n6389), .A2(n6388), .A3(n6387), .A4(n6386), .ZN(n6405) );
  AOI22D0 U2508 ( .A1(n6923), .A2(\mem[162][2] ), .B1(n6680), .B2(
        \mem[159][2] ), .ZN(n6393) );
  AOI22D0 U2509 ( .A1(n6991), .A2(\mem[148][2] ), .B1(n6659), .B2(
        \mem[181][2] ), .ZN(n6392) );
  AOI22D0 U2510 ( .A1(n6989), .A2(\mem[134][2] ), .B1(n6925), .B2(
        \mem[173][2] ), .ZN(n6391) );
  AOI22D0 U2511 ( .A1(n6814), .A2(\mem[129][2] ), .B1(n6491), .B2(
        \mem[179][2] ), .ZN(n6390) );
  ND4D0 U2512 ( .A1(n6393), .A2(n6392), .A3(n6391), .A4(n6390), .ZN(n6404) );
  AOI22D0 U2513 ( .A1(n6924), .A2(\mem[160][2] ), .B1(n6871), .B2(
        \mem[185][2] ), .ZN(n6396) );
  AOI22D0 U2514 ( .A1(n6914), .A2(\mem[133][2] ), .B1(n6922), .B2(
        \mem[157][2] ), .ZN(n6395) );
  AOI22D0 U2515 ( .A1(n6979), .A2(\mem[142][2] ), .B1(n6952), .B2(
        \mem[150][2] ), .ZN(n6394) );
  ND4D0 U2516 ( .A1(n6397), .A2(n6396), .A3(n6395), .A4(n6394), .ZN(n6403) );
  AOI22D0 U2517 ( .A1(n6880), .A2(\mem[139][2] ), .B1(n6563), .B2(
        \mem[136][2] ), .ZN(n6401) );
  AOI22D0 U2518 ( .A1(n6861), .A2(\mem[132][2] ), .B1(n6869), .B2(
        \mem[177][2] ), .ZN(n6400) );
  AOI22D0 U2519 ( .A1(n6863), .A2(\mem[183][2] ), .B1(n6964), .B2(
        \mem[158][2] ), .ZN(n6399) );
  AOI22D0 U2520 ( .A1(n6959), .A2(\mem[131][2] ), .B1(n6542), .B2(
        \mem[146][2] ), .ZN(n6398) );
  ND4D0 U2521 ( .A1(n6401), .A2(n6400), .A3(n6399), .A4(n6398), .ZN(n6402) );
  NR4D0 U2522 ( .A1(n6405), .A2(n6404), .A3(n6403), .A4(n6402), .ZN(n6427) );
  AOI22D0 U2523 ( .A1(n6901), .A2(\mem[137][2] ), .B1(n6847), .B2(
        \mem[153][2] ), .ZN(n6409) );
  AOI22D0 U2524 ( .A1(n6953), .A2(\mem[175][2] ), .B1(n6965), .B2(
        \mem[141][2] ), .ZN(n6408) );
  AOI22D0 U2525 ( .A1(n6784), .A2(\mem[156][2] ), .B1(n6733), .B2(
        \mem[186][2] ), .ZN(n6407) );
  AOI22D0 U2526 ( .A1(n6905), .A2(\mem[187][2] ), .B1(n6956), .B2(
        \mem[168][2] ), .ZN(n6406) );
  ND4D0 U2527 ( .A1(n6409), .A2(n6408), .A3(n6407), .A4(n6406), .ZN(n6425) );
  AOI22D0 U2528 ( .A1(n6967), .A2(\mem[167][2] ), .B1(n6728), .B2(
        \mem[180][2] ), .ZN(n6413) );
  AOI22D0 U2529 ( .A1(n6892), .A2(\mem[172][2] ), .B1(n6954), .B2(
        \mem[138][2] ), .ZN(n6412) );
  AOI22D0 U2530 ( .A1(n6955), .A2(\mem[149][2] ), .B1(n6995), .B2(
        \mem[151][2] ), .ZN(n6411) );
  ND4D0 U2531 ( .A1(n6413), .A2(n6412), .A3(n6411), .A4(n6410), .ZN(n6424) );
  AOI22D0 U2532 ( .A1(n6980), .A2(\mem[189][2] ), .B1(n6933), .B2(
        \mem[161][2] ), .ZN(n6417) );
  AOI22D0 U2533 ( .A1(n6890), .A2(\mem[164][2] ), .B1(n6906), .B2(
        \mem[140][2] ), .ZN(n6416) );
  AOI22D0 U2534 ( .A1(n6860), .A2(\mem[163][2] ), .B1(n6988), .B2(
        \mem[191][2] ), .ZN(n6415) );
  AOI22D0 U2535 ( .A1(n6968), .A2(\mem[169][2] ), .B1(n6992), .B2(
        \mem[182][2] ), .ZN(n6414) );
  ND4D0 U2536 ( .A1(n6417), .A2(n6416), .A3(n6415), .A4(n6414), .ZN(n6423) );
  AOI22D0 U2537 ( .A1(n6928), .A2(\mem[135][2] ), .B1(n6981), .B2(
        \mem[188][2] ), .ZN(n6421) );
  AOI22D0 U2538 ( .A1(n6934), .A2(\mem[152][2] ), .B1(n6913), .B2(
        \mem[155][2] ), .ZN(n6420) );
  AOI22D0 U2539 ( .A1(n6888), .A2(\mem[128][2] ), .B1(n6904), .B2(
        \mem[147][2] ), .ZN(n6419) );
  AOI22D0 U2540 ( .A1(n6917), .A2(\mem[174][2] ), .B1(n6982), .B2(
        \mem[130][2] ), .ZN(n6418) );
  NR4D0 U2541 ( .A1(n6425), .A2(n6424), .A3(n6423), .A4(n6422), .ZN(n6426) );
  CKND2D0 U2542 ( .A1(n6427), .A2(n6426), .ZN(n6516) );
  AOI22D0 U2543 ( .A1(n6905), .A2(\mem[123][2] ), .B1(n6804), .B2(\mem[83][2] ), .ZN(n6431) );
  AOI22D0 U2544 ( .A1(n6917), .A2(\mem[110][2] ), .B1(n6880), .B2(\mem[75][2] ), .ZN(n6430) );
  AOI22D0 U2545 ( .A1(n6861), .A2(\mem[68][2] ), .B1(n6859), .B2(\mem[116][2] ), .ZN(n6429) );
  AOI22D0 U2546 ( .A1(n6868), .A2(\mem[107][2] ), .B1(n6873), .B2(\mem[94][2] ), .ZN(n6428) );
  ND4D0 U2547 ( .A1(n6431), .A2(n6430), .A3(n6429), .A4(n6428), .ZN(n6447) );
  AOI22D0 U2548 ( .A1(n6994), .A2(\mem[126][2] ), .B1(n6862), .B2(
        \mem[104][2] ), .ZN(n6435) );
  AOI22D0 U2549 ( .A1(n6982), .A2(\mem[66][2] ), .B1(n6869), .B2(\mem[113][2] ), .ZN(n6434) );
  AOI22D0 U2550 ( .A1(n6913), .A2(\mem[91][2] ), .B1(n6791), .B2(\mem[96][2] ), 
        .ZN(n6432) );
  ND4D0 U2551 ( .A1(n6435), .A2(n6434), .A3(n6433), .A4(n6432), .ZN(n6446) );
  AOI22D0 U2552 ( .A1(n6971), .A2(\mem[102][2] ), .B1(n6871), .B2(
        \mem[121][2] ), .ZN(n6439) );
  AOI22D0 U2553 ( .A1(n6993), .A2(\mem[117][2] ), .B1(n6936), .B2(\mem[81][2] ), .ZN(n6438) );
  AOI22D0 U2554 ( .A1(n6879), .A2(\mem[122][2] ), .B1(n6658), .B2(
        \mem[114][2] ), .ZN(n6437) );
  AOI22D0 U2555 ( .A1(n6970), .A2(\mem[80][2] ), .B1(n6915), .B2(\mem[77][2] ), 
        .ZN(n6436) );
  ND4D0 U2556 ( .A1(n6439), .A2(n6438), .A3(n6437), .A4(n6436), .ZN(n6445) );
  AOI22D0 U2557 ( .A1(n6870), .A2(\mem[124][2] ), .B1(n6889), .B2(\mem[92][2] ), .ZN(n6443) );
  AOI22D0 U2558 ( .A1(n6969), .A2(\mem[82][2] ), .B1(n6901), .B2(\mem[73][2] ), 
        .ZN(n6442) );
  AOI22D0 U2559 ( .A1(n6980), .A2(\mem[125][2] ), .B1(n6882), .B2(\mem[79][2] ), .ZN(n6441) );
  AOI22D0 U2560 ( .A1(n6874), .A2(\mem[106][2] ), .B1(n6760), .B2(
        \mem[109][2] ), .ZN(n6440) );
  ND4D0 U2561 ( .A1(n6443), .A2(n6442), .A3(n6441), .A4(n6440), .ZN(n6444) );
  NR4D0 U2562 ( .A1(n6447), .A2(n6446), .A3(n6445), .A4(n6444), .ZN(n6470) );
  AOI22D0 U2563 ( .A1(n6928), .A2(\mem[71][2] ), .B1(n6891), .B2(\mem[90][2] ), 
        .ZN(n6452) );
  AOI22D0 U2564 ( .A1(n6979), .A2(\mem[78][2] ), .B1(n6902), .B2(\mem[101][2] ), .ZN(n6451) );
  AOI22D0 U2565 ( .A1(n6448), .A2(\mem[64][2] ), .B1(n6992), .B2(\mem[118][2] ), .ZN(n6450) );
  AOI22D0 U2566 ( .A1(n6976), .A2(\mem[98][2] ), .B1(n6491), .B2(\mem[115][2] ), .ZN(n6449) );
  ND4D0 U2567 ( .A1(n6452), .A2(n6451), .A3(n6450), .A4(n6449), .ZN(n6468) );
  AOI22D0 U2568 ( .A1(n6892), .A2(\mem[108][2] ), .B1(n6955), .B2(\mem[85][2] ), .ZN(n6456) );
  AOI22D0 U2569 ( .A1(n6952), .A2(\mem[86][2] ), .B1(n6863), .B2(\mem[119][2] ), .ZN(n6454) );
  AOI22D0 U2570 ( .A1(n6707), .A2(\mem[87][2] ), .B1(n6935), .B2(\mem[127][2] ), .ZN(n6453) );
  ND4D0 U2571 ( .A1(n6456), .A2(n6455), .A3(n6454), .A4(n6453), .ZN(n6467) );
  AOI22D0 U2572 ( .A1(n6883), .A2(\mem[112][2] ), .B1(n6967), .B2(
        \mem[103][2] ), .ZN(n6460) );
  AOI22D0 U2573 ( .A1(n6959), .A2(\mem[67][2] ), .B1(n6968), .B2(\mem[105][2] ), .ZN(n6459) );
  AOI22D0 U2574 ( .A1(n6927), .A2(\mem[89][2] ), .B1(n6954), .B2(\mem[74][2] ), 
        .ZN(n6458) );
  AOI22D0 U2575 ( .A1(n6953), .A2(\mem[111][2] ), .B1(n6802), .B2(\mem[88][2] ), .ZN(n6457) );
  ND4D0 U2576 ( .A1(n6460), .A2(n6459), .A3(n6458), .A4(n6457), .ZN(n6466) );
  AOI22D0 U2577 ( .A1(n6991), .A2(\mem[84][2] ), .B1(n6990), .B2(\mem[76][2] ), 
        .ZN(n6464) );
  AOI22D0 U2578 ( .A1(n6926), .A2(\mem[65][2] ), .B1(n6922), .B2(\mem[93][2] ), 
        .ZN(n6463) );
  AOI22D0 U2579 ( .A1(n6914), .A2(\mem[69][2] ), .B1(n6680), .B2(\mem[95][2] ), 
        .ZN(n6462) );
  AOI22D0 U2580 ( .A1(n6860), .A2(\mem[99][2] ), .B1(n6563), .B2(\mem[72][2] ), 
        .ZN(n6461) );
  ND4D0 U2581 ( .A1(n6464), .A2(n6463), .A3(n6462), .A4(n6461), .ZN(n6465) );
  NR4D0 U2582 ( .A1(n6468), .A2(n6467), .A3(n6466), .A4(n6465), .ZN(n6469) );
  AOI21D0 U2583 ( .A1(n6470), .A2(n6469), .B(n7004), .ZN(n6515) );
  AOI22D0 U2584 ( .A1(n6802), .A2(\mem[216][2] ), .B1(n6879), .B2(
        \mem[250][2] ), .ZN(n6474) );
  AOI22D0 U2585 ( .A1(n6614), .A2(\mem[214][2] ), .B1(n6842), .B2(
        \mem[218][2] ), .ZN(n6473) );
  AOI22D0 U2586 ( .A1(n6968), .A2(\mem[233][2] ), .B1(n6738), .B2(
        \mem[229][2] ), .ZN(n6472) );
  AOI22D0 U2587 ( .A1(n6525), .A2(\mem[227][2] ), .B1(n6933), .B2(
        \mem[225][2] ), .ZN(n6471) );
  ND4D0 U2588 ( .A1(n6474), .A2(n6473), .A3(n6472), .A4(n6471), .ZN(n6490) );
  AOI22D0 U2589 ( .A1(n6970), .A2(\mem[208][2] ), .B1(n6659), .B2(
        \mem[245][2] ), .ZN(n6477) );
  AOI22D0 U2590 ( .A1(n6953), .A2(\mem[239][2] ), .B1(n6863), .B2(
        \mem[247][2] ), .ZN(n6476) );
  AOI22D0 U2591 ( .A1(n6917), .A2(\mem[238][2] ), .B1(n6542), .B2(
        \mem[210][2] ), .ZN(n6475) );
  ND4D0 U2592 ( .A1(n6478), .A2(n6477), .A3(n6476), .A4(n6475), .ZN(n6489) );
  AOI22D0 U2593 ( .A1(n6989), .A2(\mem[198][2] ), .B1(n6837), .B2(
        \mem[207][2] ), .ZN(n6482) );
  AOI22D0 U2594 ( .A1(n6773), .A2(\mem[228][2] ), .B1(n6880), .B2(
        \mem[203][2] ), .ZN(n6481) );
  AOI22D0 U2595 ( .A1(n6925), .A2(\mem[237][2] ), .B1(n6563), .B2(
        \mem[200][2] ), .ZN(n6480) );
  AOI22D0 U2596 ( .A1(n6728), .A2(\mem[244][2] ), .B1(n6958), .B2(
        \mem[209][2] ), .ZN(n6479) );
  ND4D0 U2597 ( .A1(n6482), .A2(n6481), .A3(n6480), .A4(n6479), .ZN(n6488) );
  AOI22D0 U2598 ( .A1(n6959), .A2(\mem[195][2] ), .B1(n6868), .B2(
        \mem[235][2] ), .ZN(n6486) );
  AOI22D0 U2599 ( .A1(n6814), .A2(\mem[193][2] ), .B1(n6789), .B2(
        \mem[254][2] ), .ZN(n6485) );
  AOI22D0 U2600 ( .A1(n6680), .A2(\mem[223][2] ), .B1(n6924), .B2(
        \mem[224][2] ), .ZN(n6484) );
  AOI22D0 U2601 ( .A1(n6530), .A2(\mem[251][2] ), .B1(n6790), .B2(
        \mem[219][2] ), .ZN(n6483) );
  ND4D0 U2602 ( .A1(n6486), .A2(n6485), .A3(n6484), .A4(n6483), .ZN(n6487) );
  NR4D0 U2603 ( .A1(n6490), .A2(n6489), .A3(n6488), .A4(n6487), .ZN(n6513) );
  AOI22D0 U2604 ( .A1(n6759), .A2(\mem[206][2] ), .B1(n6992), .B2(
        \mem[246][2] ), .ZN(n6495) );
  AOI22D0 U2605 ( .A1(n6874), .A2(\mem[234][2] ), .B1(n6976), .B2(
        \mem[226][2] ), .ZN(n6494) );
  AOI22D0 U2606 ( .A1(n6928), .A2(\mem[199][2] ), .B1(n6491), .B2(
        \mem[243][2] ), .ZN(n6493) );
  ND4D0 U2607 ( .A1(n6495), .A2(n6494), .A3(n6493), .A4(n6492), .ZN(n6511) );
  AOI22D0 U2608 ( .A1(n6957), .A2(\mem[249][2] ), .B1(n6906), .B2(
        \mem[204][2] ), .ZN(n6499) );
  AOI22D0 U2609 ( .A1(n6904), .A2(\mem[211][2] ), .B1(n6774), .B2(
        \mem[241][2] ), .ZN(n6498) );
  AOI22D0 U2610 ( .A1(n6955), .A2(\mem[213][2] ), .B1(n6956), .B2(
        \mem[232][2] ), .ZN(n6497) );
  AOI22D0 U2611 ( .A1(n6914), .A2(\mem[197][2] ), .B1(n6995), .B2(
        \mem[215][2] ), .ZN(n6496) );
  ND4D0 U2612 ( .A1(n6499), .A2(n6498), .A3(n6497), .A4(n6496), .ZN(n6510) );
  AOI22D0 U2613 ( .A1(n6883), .A2(\mem[240][2] ), .B1(n6915), .B2(
        \mem[205][2] ), .ZN(n6503) );
  AOI22D0 U2614 ( .A1(n6847), .A2(\mem[217][2] ), .B1(n6954), .B2(
        \mem[202][2] ), .ZN(n6502) );
  AOI22D0 U2615 ( .A1(n6861), .A2(\mem[196][2] ), .B1(n6888), .B2(
        \mem[192][2] ), .ZN(n6501) );
  AOI22D0 U2616 ( .A1(n6658), .A2(\mem[242][2] ), .B1(n6698), .B2(
        \mem[194][2] ), .ZN(n6500) );
  AOI22D0 U2617 ( .A1(n6980), .A2(\mem[253][2] ), .B1(n6889), .B2(
        \mem[220][2] ), .ZN(n6507) );
  AOI22D0 U2618 ( .A1(n6981), .A2(\mem[252][2] ), .B1(n6964), .B2(
        \mem[222][2] ), .ZN(n6506) );
  AOI22D0 U2619 ( .A1(n6809), .A2(\mem[201][2] ), .B1(n6912), .B2(
        \mem[248][2] ), .ZN(n6505) );
  AOI22D0 U2620 ( .A1(n6892), .A2(\mem[236][2] ), .B1(n6829), .B2(
        \mem[230][2] ), .ZN(n6504) );
  ND4D0 U2621 ( .A1(n6507), .A2(n6506), .A3(n6505), .A4(n6504), .ZN(n6508) );
  NR4D0 U2622 ( .A1(n6511), .A2(n6510), .A3(n6509), .A4(n6508), .ZN(n6512) );
  AOI21D0 U2623 ( .A1(n6513), .A2(n6512), .B(n6945), .ZN(n6514) );
  AOI211D0 U2624 ( .A1(n6951), .A2(n6516), .B(n6515), .C(n6514), .ZN(n6540) );
  AOI22D0 U2625 ( .A1(n6862), .A2(\mem[40][2] ), .B1(n6912), .B2(\mem[56][2] ), 
        .ZN(n6520) );
  AOI22D0 U2626 ( .A1(n6928), .A2(\mem[7][2] ), .B1(n6957), .B2(\mem[57][2] ), 
        .ZN(n6519) );
  AOI22D0 U2627 ( .A1(n6968), .A2(\mem[41][2] ), .B1(n6882), .B2(\mem[15][2] ), 
        .ZN(n6518) );
  AOI22D0 U2628 ( .A1(n6958), .A2(\mem[17][2] ), .B1(n6836), .B2(\mem[10][2] ), 
        .ZN(n6517) );
  ND4D0 U2629 ( .A1(n6520), .A2(n6519), .A3(n6518), .A4(n6517), .ZN(n6538) );
  AOI22D0 U2630 ( .A1(n6890), .A2(\mem[36][2] ), .B1(n6926), .B2(\mem[1][2] ), 
        .ZN(n6524) );
  AOI22D0 U2631 ( .A1(n6971), .A2(\mem[38][2] ), .B1(n6658), .B2(\mem[50][2] ), 
        .ZN(n6523) );
  AOI22D0 U2632 ( .A1(n6953), .A2(\mem[47][2] ), .B1(n6965), .B2(\mem[13][2] ), 
        .ZN(n6522) );
  AOI22D0 U2633 ( .A1(n6863), .A2(\mem[55][2] ), .B1(n6859), .B2(\mem[52][2] ), 
        .ZN(n6521) );
  ND4D0 U2634 ( .A1(n6524), .A2(n6523), .A3(n6522), .A4(n6521), .ZN(n6537) );
  AOI22D0 U2635 ( .A1(n6802), .A2(\mem[24][2] ), .B1(n6933), .B2(\mem[33][2] ), 
        .ZN(n6528) );
  AOI22D0 U2636 ( .A1(n6614), .A2(\mem[22][2] ), .B1(n6869), .B2(\mem[49][2] ), 
        .ZN(n6527) );
  AOI22D0 U2637 ( .A1(n6917), .A2(\mem[46][2] ), .B1(n6888), .B2(\mem[0][2] ), 
        .ZN(n6526) );
  AOI22D0 U2638 ( .A1(n6969), .A2(\mem[18][2] ), .B1(n6698), .B2(\mem[2][2] ), 
        .ZN(n6534) );
  AOI22D0 U2639 ( .A1(n6989), .A2(\mem[6][2] ), .B1(n6563), .B2(\mem[8][2] ), 
        .ZN(n6533) );
  AOI22D0 U2640 ( .A1(n6530), .A2(\mem[59][2] ), .B1(n6967), .B2(\mem[39][2] ), 
        .ZN(n6532) );
  AOI22D0 U2641 ( .A1(n6868), .A2(\mem[43][2] ), .B1(n6790), .B2(\mem[27][2] ), 
        .ZN(n6531) );
  ND4D0 U2642 ( .A1(n6534), .A2(n6533), .A3(n6532), .A4(n6531), .ZN(n6535) );
  NR4D0 U2643 ( .A1(n6538), .A2(n6537), .A3(n6536), .A4(n6535), .ZN(n6539) );
  AOI32D0 U2644 ( .A1(n6541), .A2(n6540), .A3(n6539), .B1(n6856), .B2(n6540), 
        .ZN(dout[2]) );
  AOI22D0 U2645 ( .A1(n6814), .A2(\mem[65][3] ), .B1(n6542), .B2(\mem[82][3] ), 
        .ZN(n6546) );
  AOI22D0 U2646 ( .A1(n6924), .A2(\mem[96][3] ), .B1(n6955), .B2(\mem[85][3] ), 
        .ZN(n6545) );
  AOI22D0 U2647 ( .A1(n6873), .A2(\mem[94][3] ), .B1(n6992), .B2(\mem[118][3] ), .ZN(n6544) );
  AOI22D0 U2648 ( .A1(n6991), .A2(\mem[84][3] ), .B1(n6829), .B2(\mem[102][3] ), .ZN(n6543) );
  ND4D0 U2649 ( .A1(n6546), .A2(n6545), .A3(n6544), .A4(n6543), .ZN(n6562) );
  AOI22D0 U2650 ( .A1(n6988), .A2(\mem[127][3] ), .B1(n6760), .B2(
        \mem[109][3] ), .ZN(n6550) );
  AOI22D0 U2651 ( .A1(n6905), .A2(\mem[123][3] ), .B1(n6680), .B2(\mem[95][3] ), .ZN(n6549) );
  AOI22D0 U2652 ( .A1(n6888), .A2(\mem[64][3] ), .B1(n6913), .B2(\mem[91][3] ), 
        .ZN(n6548) );
  AOI22D0 U2653 ( .A1(n6891), .A2(\mem[90][3] ), .B1(n6836), .B2(\mem[74][3] ), 
        .ZN(n6547) );
  ND4D0 U2654 ( .A1(n6550), .A2(n6549), .A3(n6548), .A4(n6547), .ZN(n6561) );
  AOI22D0 U2655 ( .A1(n6639), .A2(\mem[103][3] ), .B1(n6828), .B2(
        \mem[120][3] ), .ZN(n6553) );
  AOI22D0 U2656 ( .A1(n6981), .A2(\mem[124][3] ), .B1(n6658), .B2(
        \mem[114][3] ), .ZN(n6552) );
  AOI22D0 U2657 ( .A1(n6970), .A2(\mem[80][3] ), .B1(n6957), .B2(\mem[121][3] ), .ZN(n6551) );
  ND4D0 U2658 ( .A1(n6554), .A2(n6553), .A3(n6552), .A4(n6551), .ZN(n6560) );
  AOI22D0 U2659 ( .A1(n6953), .A2(\mem[111][3] ), .B1(n6990), .B2(\mem[76][3] ), .ZN(n6558) );
  AOI22D0 U2660 ( .A1(n6880), .A2(\mem[75][3] ), .B1(n6804), .B2(\mem[83][3] ), 
        .ZN(n6557) );
  AOI22D0 U2661 ( .A1(n6917), .A2(\mem[110][3] ), .B1(n6847), .B2(\mem[89][3] ), .ZN(n6556) );
  AOI22D0 U2662 ( .A1(n6907), .A2(\mem[67][3] ), .B1(n6728), .B2(\mem[116][3] ), .ZN(n6555) );
  ND4D0 U2663 ( .A1(n6558), .A2(n6557), .A3(n6556), .A4(n6555), .ZN(n6559) );
  NR4D0 U2664 ( .A1(n6562), .A2(n6561), .A3(n6560), .A4(n6559), .ZN(n6722) );
  AOI22D0 U2665 ( .A1(n6905), .A2(\mem[187][3] ), .B1(n6992), .B2(
        \mem[182][3] ), .ZN(n6567) );
  AOI22D0 U2666 ( .A1(n6959), .A2(\mem[131][3] ), .B1(n6914), .B2(
        \mem[133][3] ), .ZN(n6566) );
  AOI22D0 U2667 ( .A1(n6903), .A2(\mem[179][3] ), .B1(n6994), .B2(
        \mem[190][3] ), .ZN(n6565) );
  AOI22D0 U2668 ( .A1(n6802), .A2(\mem[152][3] ), .B1(n6563), .B2(
        \mem[136][3] ), .ZN(n6564) );
  ND4D0 U2669 ( .A1(n6567), .A2(n6566), .A3(n6565), .A4(n6564), .ZN(n6583) );
  AOI22D0 U2670 ( .A1(n6863), .A2(\mem[183][3] ), .B1(n6733), .B2(
        \mem[186][3] ), .ZN(n6571) );
  AOI22D0 U2671 ( .A1(n6728), .A2(\mem[180][3] ), .B1(n6956), .B2(
        \mem[168][3] ), .ZN(n6570) );
  AOI22D0 U2672 ( .A1(n6983), .A2(\mem[176][3] ), .B1(n6933), .B2(
        \mem[161][3] ), .ZN(n6569) );
  AOI22D0 U2673 ( .A1(n6952), .A2(\mem[150][3] ), .B1(n6882), .B2(
        \mem[143][3] ), .ZN(n6568) );
  ND4D0 U2674 ( .A1(n6571), .A2(n6570), .A3(n6569), .A4(n6568), .ZN(n6582) );
  AOI22D0 U2675 ( .A1(n6928), .A2(\mem[135][3] ), .B1(n6970), .B2(
        \mem[144][3] ), .ZN(n6575) );
  AOI22D0 U2676 ( .A1(n6889), .A2(\mem[156][3] ), .B1(n6958), .B2(
        \mem[145][3] ), .ZN(n6574) );
  AOI22D0 U2677 ( .A1(n6890), .A2(\mem[164][3] ), .B1(n6912), .B2(
        \mem[184][3] ), .ZN(n6573) );
  AOI22D0 U2678 ( .A1(n6991), .A2(\mem[148][3] ), .B1(n6836), .B2(
        \mem[138][3] ), .ZN(n6572) );
  AOI22D0 U2679 ( .A1(n6926), .A2(\mem[129][3] ), .B1(n6922), .B2(
        \mem[157][3] ), .ZN(n6579) );
  AOI22D0 U2680 ( .A1(n6925), .A2(\mem[173][3] ), .B1(n6774), .B2(
        \mem[177][3] ), .ZN(n6578) );
  AOI22D0 U2681 ( .A1(n6892), .A2(\mem[172][3] ), .B1(n6659), .B2(
        \mem[181][3] ), .ZN(n6576) );
  ND4D0 U2682 ( .A1(n6579), .A2(n6578), .A3(n6577), .A4(n6576), .ZN(n6580) );
  NR4D0 U2683 ( .A1(n6583), .A2(n6582), .A3(n6581), .A4(n6580), .ZN(n6605) );
  AOI22D0 U2684 ( .A1(n6680), .A2(\mem[159][3] ), .B1(n6966), .B2(
        \mem[178][3] ), .ZN(n6587) );
  AOI22D0 U2685 ( .A1(n6935), .A2(\mem[191][3] ), .B1(n6871), .B2(
        \mem[185][3] ), .ZN(n6586) );
  AOI22D0 U2686 ( .A1(n6967), .A2(\mem[167][3] ), .B1(n6968), .B2(
        \mem[169][3] ), .ZN(n6585) );
  AOI22D0 U2687 ( .A1(n6976), .A2(\mem[162][3] ), .B1(n6847), .B2(
        \mem[153][3] ), .ZN(n6584) );
  ND4D0 U2688 ( .A1(n6587), .A2(n6586), .A3(n6585), .A4(n6584), .ZN(n6603) );
  AOI22D0 U2689 ( .A1(n6969), .A2(\mem[146][3] ), .B1(n6915), .B2(
        \mem[141][3] ), .ZN(n6591) );
  AOI22D0 U2690 ( .A1(n6981), .A2(\mem[188][3] ), .B1(n6888), .B2(
        \mem[128][3] ), .ZN(n6590) );
  AOI22D0 U2691 ( .A1(n6980), .A2(\mem[189][3] ), .B1(n6829), .B2(
        \mem[166][3] ), .ZN(n6589) );
  AOI22D0 U2692 ( .A1(n6989), .A2(\mem[134][3] ), .B1(n6902), .B2(
        \mem[165][3] ), .ZN(n6588) );
  ND4D0 U2693 ( .A1(n6591), .A2(n6590), .A3(n6589), .A4(n6588), .ZN(n6602) );
  AOI22D0 U2694 ( .A1(n6809), .A2(\mem[137][3] ), .B1(n6707), .B2(
        \mem[151][3] ), .ZN(n6595) );
  AOI22D0 U2695 ( .A1(n6749), .A2(\mem[171][3] ), .B1(n6874), .B2(
        \mem[170][3] ), .ZN(n6594) );
  AOI22D0 U2696 ( .A1(n6982), .A2(\mem[130][3] ), .B1(n6873), .B2(
        \mem[158][3] ), .ZN(n6593) );
  AOI22D0 U2697 ( .A1(n6953), .A2(\mem[175][3] ), .B1(n6835), .B2(
        \mem[132][3] ), .ZN(n6592) );
  ND4D0 U2698 ( .A1(n6595), .A2(n6594), .A3(n6593), .A4(n6592), .ZN(n6601) );
  AOI22D0 U2699 ( .A1(n6924), .A2(\mem[160][3] ), .B1(n6904), .B2(
        \mem[147][3] ), .ZN(n6599) );
  AOI22D0 U2700 ( .A1(n6860), .A2(\mem[163][3] ), .B1(n6916), .B2(
        \mem[149][3] ), .ZN(n6597) );
  AOI22D0 U2701 ( .A1(n6979), .A2(\mem[142][3] ), .B1(n6891), .B2(
        \mem[154][3] ), .ZN(n6596) );
  ND4D0 U2702 ( .A1(n6599), .A2(n6598), .A3(n6597), .A4(n6596), .ZN(n6600) );
  NR4D0 U2703 ( .A1(n6603), .A2(n6602), .A3(n6601), .A4(n6600), .ZN(n6604) );
  CKND2D0 U2704 ( .A1(n6605), .A2(n6604), .ZN(n6697) );
  AOI22D0 U2705 ( .A1(n6959), .A2(\mem[3][3] ), .B1(n6979), .B2(\mem[14][3] ), 
        .ZN(n6609) );
  AOI22D0 U2706 ( .A1(n6924), .A2(\mem[32][3] ), .B1(n6837), .B2(\mem[15][3] ), 
        .ZN(n6608) );
  AOI22D0 U2707 ( .A1(n6879), .A2(\mem[58][3] ), .B1(n6976), .B2(\mem[34][3] ), 
        .ZN(n6607) );
  AOI22D0 U2708 ( .A1(n6728), .A2(\mem[52][3] ), .B1(n6992), .B2(\mem[54][3] ), 
        .ZN(n6606) );
  ND4D0 U2709 ( .A1(n6609), .A2(n6608), .A3(n6607), .A4(n6606), .ZN(n6626) );
  AOI22D0 U2710 ( .A1(n6980), .A2(\mem[61][3] ), .B1(n6957), .B2(\mem[57][3] ), 
        .ZN(n6613) );
  AOI22D0 U2711 ( .A1(n6969), .A2(\mem[18][3] ), .B1(n6738), .B2(\mem[37][3] ), 
        .ZN(n6612) );
  AOI22D0 U2712 ( .A1(n6790), .A2(\mem[27][3] ), .B1(n6978), .B2(\mem[8][3] ), 
        .ZN(n6611) );
  AOI22D0 U2713 ( .A1(n6890), .A2(\mem[36][3] ), .B1(n6956), .B2(\mem[40][3] ), 
        .ZN(n6610) );
  ND4D0 U2714 ( .A1(n6613), .A2(n6612), .A3(n6611), .A4(n6610), .ZN(n6625) );
  AOI22D0 U2715 ( .A1(n6970), .A2(\mem[16][3] ), .B1(n6658), .B2(\mem[50][3] ), 
        .ZN(n6618) );
  AOI22D0 U2716 ( .A1(n6971), .A2(\mem[38][3] ), .B1(n6912), .B2(\mem[56][3] ), 
        .ZN(n6617) );
  AOI22D0 U2717 ( .A1(n6614), .A2(\mem[22][3] ), .B1(n6922), .B2(\mem[29][3] ), 
        .ZN(n6616) );
  AOI22D0 U2718 ( .A1(n6880), .A2(\mem[11][3] ), .B1(n6903), .B2(\mem[51][3] ), 
        .ZN(n6615) );
  ND4D0 U2719 ( .A1(n6618), .A2(n6617), .A3(n6616), .A4(n6615), .ZN(n6624) );
  AOI22D0 U2720 ( .A1(n6860), .A2(\mem[35][3] ), .B1(n6994), .B2(\mem[62][3] ), 
        .ZN(n6621) );
  AOI22D0 U2721 ( .A1(n6680), .A2(\mem[31][3] ), .B1(n6904), .B2(\mem[19][3] ), 
        .ZN(n6620) );
  AOI22D0 U2722 ( .A1(n6803), .A2(\mem[55][3] ), .B1(n6935), .B2(\mem[63][3] ), 
        .ZN(n6619) );
  ND4D0 U2723 ( .A1(n6622), .A2(n6621), .A3(n6620), .A4(n6619), .ZN(n6623) );
  NR4D0 U2724 ( .A1(n6626), .A2(n6625), .A3(n6624), .A4(n6623), .ZN(n6649) );
  AOI22D0 U2725 ( .A1(n6928), .A2(\mem[7][3] ), .B1(n6968), .B2(\mem[41][3] ), 
        .ZN(n6630) );
  AOI22D0 U2726 ( .A1(n6953), .A2(\mem[47][3] ), .B1(n6883), .B2(\mem[48][3] ), 
        .ZN(n6629) );
  AOI22D0 U2727 ( .A1(n6989), .A2(\mem[6][3] ), .B1(n6933), .B2(\mem[33][3] ), 
        .ZN(n6628) );
  AOI22D0 U2728 ( .A1(n6916), .A2(\mem[21][3] ), .B1(n6873), .B2(\mem[30][3] ), 
        .ZN(n6627) );
  ND4D0 U2729 ( .A1(n6630), .A2(n6629), .A3(n6628), .A4(n6627), .ZN(n6647) );
  AOI22D0 U2730 ( .A1(n6874), .A2(\mem[42][3] ), .B1(n6760), .B2(\mem[45][3] ), 
        .ZN(n6634) );
  AOI22D0 U2731 ( .A1(n6954), .A2(\mem[10][3] ), .B1(n6990), .B2(\mem[12][3] ), 
        .ZN(n6633) );
  AOI22D0 U2732 ( .A1(n6905), .A2(\mem[59][3] ), .B1(n6926), .B2(\mem[1][3] ), 
        .ZN(n6632) );
  AOI22D0 U2733 ( .A1(n6917), .A2(\mem[46][3] ), .B1(n6659), .B2(\mem[53][3] ), 
        .ZN(n6631) );
  ND4D0 U2734 ( .A1(n6634), .A2(n6633), .A3(n6632), .A4(n6631), .ZN(n6646) );
  AOI22D0 U2735 ( .A1(n6870), .A2(\mem[60][3] ), .B1(n6835), .B2(\mem[4][3] ), 
        .ZN(n6638) );
  AOI22D0 U2736 ( .A1(n6707), .A2(\mem[23][3] ), .B1(n6965), .B2(\mem[13][3] ), 
        .ZN(n6637) );
  AOI22D0 U2737 ( .A1(n6914), .A2(\mem[5][3] ), .B1(n6901), .B2(\mem[9][3] ), 
        .ZN(n6636) );
  ND4D0 U2738 ( .A1(n6638), .A2(n6637), .A3(n6636), .A4(n6635), .ZN(n6645) );
  AOI22D0 U2739 ( .A1(n6991), .A2(\mem[20][3] ), .B1(n6888), .B2(\mem[0][3] ), 
        .ZN(n6643) );
  AOI22D0 U2740 ( .A1(n6892), .A2(\mem[44][3] ), .B1(n6842), .B2(\mem[26][3] ), 
        .ZN(n6642) );
  AOI22D0 U2741 ( .A1(n6749), .A2(\mem[43][3] ), .B1(n6639), .B2(\mem[39][3] ), 
        .ZN(n6641) );
  AOI22D0 U2742 ( .A1(n6934), .A2(\mem[24][3] ), .B1(n6958), .B2(\mem[17][3] ), 
        .ZN(n6640) );
  ND4D0 U2743 ( .A1(n6643), .A2(n6642), .A3(n6641), .A4(n6640), .ZN(n6644) );
  NR4D0 U2744 ( .A1(n6647), .A2(n6646), .A3(n6645), .A4(n6644), .ZN(n6648) );
  AOI22D0 U2745 ( .A1(n6959), .A2(\mem[195][3] ), .B1(n6979), .B2(
        \mem[206][3] ), .ZN(n6653) );
  AOI22D0 U2746 ( .A1(n6913), .A2(\mem[219][3] ), .B1(n6873), .B2(
        \mem[222][3] ), .ZN(n6652) );
  AOI22D0 U2747 ( .A1(n6905), .A2(\mem[251][3] ), .B1(n6698), .B2(
        \mem[194][3] ), .ZN(n6651) );
  AOI22D0 U2748 ( .A1(n6969), .A2(\mem[210][3] ), .B1(n6990), .B2(
        \mem[204][3] ), .ZN(n6650) );
  ND4D0 U2749 ( .A1(n6653), .A2(n6652), .A3(n6651), .A4(n6650), .ZN(n6671) );
  AOI22D0 U2750 ( .A1(n6967), .A2(\mem[231][3] ), .B1(n6863), .B2(
        \mem[247][3] ), .ZN(n6657) );
  AOI22D0 U2751 ( .A1(n6980), .A2(\mem[253][3] ), .B1(n6881), .B2(
        \mem[208][3] ), .ZN(n6656) );
  AOI22D0 U2752 ( .A1(n6883), .A2(\mem[240][3] ), .B1(n6859), .B2(
        \mem[244][3] ), .ZN(n6655) );
  AOI22D0 U2753 ( .A1(n6917), .A2(\mem[238][3] ), .B1(n6928), .B2(
        \mem[199][3] ), .ZN(n6654) );
  AOI22D0 U2754 ( .A1(n6870), .A2(\mem[252][3] ), .B1(n6658), .B2(
        \mem[242][3] ), .ZN(n6663) );
  AOI22D0 U2755 ( .A1(n6879), .A2(\mem[250][3] ), .B1(n6659), .B2(
        \mem[245][3] ), .ZN(n6662) );
  AOI22D0 U2756 ( .A1(n6991), .A2(\mem[212][3] ), .B1(n6791), .B2(
        \mem[224][3] ), .ZN(n6660) );
  ND4D0 U2757 ( .A1(n6663), .A2(n6662), .A3(n6661), .A4(n6660), .ZN(n6669) );
  AOI22D0 U2758 ( .A1(n6892), .A2(\mem[236][3] ), .B1(n6923), .B2(
        \mem[226][3] ), .ZN(n6667) );
  AOI22D0 U2759 ( .A1(n6868), .A2(\mem[235][3] ), .B1(n6989), .B2(
        \mem[198][3] ), .ZN(n6666) );
  AOI22D0 U2760 ( .A1(n6837), .A2(\mem[207][3] ), .B1(n6828), .B2(
        \mem[248][3] ), .ZN(n6665) );
  AOI22D0 U2761 ( .A1(n6933), .A2(\mem[225][3] ), .B1(n6707), .B2(
        \mem[215][3] ), .ZN(n6664) );
  ND4D0 U2762 ( .A1(n6667), .A2(n6666), .A3(n6665), .A4(n6664), .ZN(n6668) );
  NR4D0 U2763 ( .A1(n6671), .A2(n6670), .A3(n6669), .A4(n6668), .ZN(n6694) );
  AOI22D0 U2764 ( .A1(n6754), .A2(\mem[197][3] ), .B1(n6862), .B2(
        \mem[232][3] ), .ZN(n6675) );
  AOI22D0 U2765 ( .A1(n6842), .A2(\mem[218][3] ), .B1(n6902), .B2(
        \mem[229][3] ), .ZN(n6674) );
  AOI22D0 U2766 ( .A1(n6874), .A2(\mem[234][3] ), .B1(n6922), .B2(
        \mem[221][3] ), .ZN(n6673) );
  AOI22D0 U2767 ( .A1(n6802), .A2(\mem[216][3] ), .B1(n6957), .B2(
        \mem[249][3] ), .ZN(n6672) );
  ND4D0 U2768 ( .A1(n6675), .A2(n6674), .A3(n6673), .A4(n6672), .ZN(n6692) );
  AOI22D0 U2769 ( .A1(n6927), .A2(\mem[217][3] ), .B1(n6954), .B2(
        \mem[202][3] ), .ZN(n6679) );
  AOI22D0 U2770 ( .A1(n6926), .A2(\mem[193][3] ), .B1(n6903), .B2(
        \mem[243][3] ), .ZN(n6678) );
  AOI22D0 U2771 ( .A1(n6953), .A2(\mem[239][3] ), .B1(n6869), .B2(
        \mem[241][3] ), .ZN(n6677) );
  AOI22D0 U2772 ( .A1(n6880), .A2(\mem[203][3] ), .B1(n6888), .B2(
        \mem[192][3] ), .ZN(n6676) );
  ND4D0 U2773 ( .A1(n6679), .A2(n6678), .A3(n6677), .A4(n6676), .ZN(n6691) );
  AOI22D0 U2774 ( .A1(n6968), .A2(\mem[233][3] ), .B1(n6915), .B2(
        \mem[205][3] ), .ZN(n6684) );
  AOI22D0 U2775 ( .A1(n6952), .A2(\mem[214][3] ), .B1(n6680), .B2(
        \mem[223][3] ), .ZN(n6682) );
  AOI22D0 U2776 ( .A1(n6901), .A2(\mem[201][3] ), .B1(n6978), .B2(
        \mem[200][3] ), .ZN(n6681) );
  ND4D0 U2777 ( .A1(n6684), .A2(n6683), .A3(n6682), .A4(n6681), .ZN(n6690) );
  AOI22D0 U2778 ( .A1(n6971), .A2(\mem[230][3] ), .B1(n6904), .B2(
        \mem[211][3] ), .ZN(n6688) );
  AOI22D0 U2779 ( .A1(n6988), .A2(\mem[255][3] ), .B1(n6992), .B2(
        \mem[246][3] ), .ZN(n6687) );
  AOI22D0 U2780 ( .A1(n6861), .A2(\mem[196][3] ), .B1(n6958), .B2(
        \mem[209][3] ), .ZN(n6686) );
  AOI22D0 U2781 ( .A1(n6784), .A2(\mem[220][3] ), .B1(n6955), .B2(
        \mem[213][3] ), .ZN(n6685) );
  ND4D0 U2782 ( .A1(n6688), .A2(n6687), .A3(n6686), .A4(n6685), .ZN(n6689) );
  NR4D0 U2783 ( .A1(n6692), .A2(n6691), .A3(n6690), .A4(n6689), .ZN(n6693) );
  AOI21D0 U2784 ( .A1(n6694), .A2(n6693), .B(n6945), .ZN(n6695) );
  AOI211D0 U2785 ( .A1(n6951), .A2(n6697), .B(n6696), .C(n6695), .ZN(n6721) );
  AOI22D0 U2786 ( .A1(n6993), .A2(\mem[117][3] ), .B1(n6698), .B2(\mem[66][3] ), .ZN(n6702) );
  AOI22D0 U2787 ( .A1(n6989), .A2(\mem[70][3] ), .B1(n6902), .B2(\mem[101][3] ), .ZN(n6700) );
  AOI22D0 U2788 ( .A1(n6914), .A2(\mem[69][3] ), .B1(n6874), .B2(\mem[106][3] ), .ZN(n6699) );
  ND4D0 U2789 ( .A1(n6702), .A2(n6701), .A3(n6700), .A4(n6699), .ZN(n6719) );
  AOI22D0 U2790 ( .A1(n6868), .A2(\mem[107][3] ), .B1(n6933), .B2(\mem[97][3] ), .ZN(n6706) );
  AOI22D0 U2791 ( .A1(n6903), .A2(\mem[115][3] ), .B1(n6774), .B2(
        \mem[113][3] ), .ZN(n6705) );
  AOI22D0 U2792 ( .A1(n6860), .A2(\mem[99][3] ), .B1(n6879), .B2(\mem[122][3] ), .ZN(n6704) );
  AOI22D0 U2793 ( .A1(n6802), .A2(\mem[88][3] ), .B1(n6901), .B2(\mem[73][3] ), 
        .ZN(n6703) );
  ND4D0 U2794 ( .A1(n6706), .A2(n6705), .A3(n6704), .A4(n6703), .ZN(n6718) );
  AOI22D0 U2795 ( .A1(n6861), .A2(\mem[68][3] ), .B1(n6958), .B2(\mem[81][3] ), 
        .ZN(n6711) );
  AOI22D0 U2796 ( .A1(n6979), .A2(\mem[78][3] ), .B1(n6882), .B2(\mem[79][3] ), 
        .ZN(n6710) );
  AOI22D0 U2797 ( .A1(n6928), .A2(\mem[71][3] ), .B1(n6956), .B2(\mem[104][3] ), .ZN(n6709) );
  AOI22D0 U2798 ( .A1(n6980), .A2(\mem[125][3] ), .B1(n6707), .B2(\mem[87][3] ), .ZN(n6708) );
  ND4D0 U2799 ( .A1(n6711), .A2(n6710), .A3(n6709), .A4(n6708), .ZN(n6717) );
  AOI22D0 U2800 ( .A1(n6983), .A2(\mem[112][3] ), .B1(n6863), .B2(
        \mem[119][3] ), .ZN(n6715) );
  AOI22D0 U2801 ( .A1(n6994), .A2(\mem[126][3] ), .B1(n6965), .B2(\mem[77][3] ), .ZN(n6714) );
  AOI22D0 U2802 ( .A1(n6923), .A2(\mem[98][3] ), .B1(n6978), .B2(\mem[72][3] ), 
        .ZN(n6713) );
  AOI22D0 U2803 ( .A1(n6890), .A2(\mem[100][3] ), .B1(n6968), .B2(
        \mem[105][3] ), .ZN(n6712) );
  ND4D0 U2804 ( .A1(n6715), .A2(n6714), .A3(n6713), .A4(n6712), .ZN(n6716) );
  NR4D0 U2805 ( .A1(n6719), .A2(n6718), .A3(n6717), .A4(n6716), .ZN(n6720) );
  AOI22D0 U2806 ( .A1(n6847), .A2(\mem[89][1] ), .B1(n6904), .B2(\mem[83][1] ), 
        .ZN(n6726) );
  AOI22D0 U2807 ( .A1(n6775), .A2(\mem[108][1] ), .B1(n6784), .B2(\mem[92][1] ), .ZN(n6725) );
  AOI22D0 U2808 ( .A1(n6905), .A2(\mem[123][1] ), .B1(n6901), .B2(\mem[73][1] ), .ZN(n6724) );
  AOI22D0 U2809 ( .A1(n6922), .A2(\mem[93][1] ), .B1(n6882), .B2(\mem[79][1] ), 
        .ZN(n6723) );
  ND4D0 U2810 ( .A1(n6726), .A2(n6725), .A3(n6724), .A4(n6723), .ZN(n6746) );
  AOI22D0 U2811 ( .A1(n6934), .A2(\mem[88][1] ), .B1(n6903), .B2(\mem[115][1] ), .ZN(n6732) );
  AOI22D0 U2812 ( .A1(n6727), .A2(\mem[106][1] ), .B1(n6680), .B2(\mem[95][1] ), .ZN(n6731) );
  AOI22D0 U2813 ( .A1(n6749), .A2(\mem[107][1] ), .B1(n6924), .B2(\mem[96][1] ), .ZN(n6730) );
  AOI22D0 U2814 ( .A1(n6728), .A2(\mem[116][1] ), .B1(n6760), .B2(
        \mem[109][1] ), .ZN(n6729) );
  ND4D0 U2815 ( .A1(n6732), .A2(n6731), .A3(n6730), .A4(n6729), .ZN(n6745) );
  AOI22D0 U2816 ( .A1(n6888), .A2(\mem[64][1] ), .B1(n6733), .B2(\mem[122][1] ), .ZN(n6737) );
  AOI22D0 U2817 ( .A1(n6814), .A2(\mem[65][1] ), .B1(n6861), .B2(\mem[68][1] ), 
        .ZN(n6736) );
  AOI22D0 U2818 ( .A1(n6890), .A2(\mem[100][1] ), .B1(n6863), .B2(
        \mem[119][1] ), .ZN(n6735) );
  AOI22D0 U2819 ( .A1(n6928), .A2(\mem[71][1] ), .B1(n6754), .B2(\mem[69][1] ), 
        .ZN(n6734) );
  ND4D0 U2820 ( .A1(n6737), .A2(n6736), .A3(n6735), .A4(n6734), .ZN(n6744) );
  AOI22D0 U2821 ( .A1(n6913), .A2(\mem[91][1] ), .B1(n6828), .B2(\mem[120][1] ), .ZN(n6742) );
  AOI22D0 U2822 ( .A1(n6917), .A2(\mem[110][1] ), .B1(n6880), .B2(\mem[75][1] ), .ZN(n6740) );
  AOI22D0 U2823 ( .A1(n6891), .A2(\mem[90][1] ), .B1(n6738), .B2(\mem[101][1] ), .ZN(n6739) );
  ND4D0 U2824 ( .A1(n6742), .A2(n6741), .A3(n6740), .A4(n6739), .ZN(n6743) );
  NR4D0 U2825 ( .A1(n6746), .A2(n6745), .A3(n6744), .A4(n6743), .ZN(n7007) );
  AOI22D0 U2826 ( .A1(n6747), .A2(\mem[148][1] ), .B1(n6978), .B2(
        \mem[136][1] ), .ZN(n6753) );
  AOI22D0 U2827 ( .A1(n6861), .A2(\mem[132][1] ), .B1(n6879), .B2(
        \mem[186][1] ), .ZN(n6752) );
  AOI22D0 U2828 ( .A1(n6830), .A2(\mem[135][1] ), .B1(n6748), .B2(
        \mem[169][1] ), .ZN(n6751) );
  AOI22D0 U2829 ( .A1(n6749), .A2(\mem[171][1] ), .B1(n6903), .B2(
        \mem[179][1] ), .ZN(n6750) );
  ND4D0 U2830 ( .A1(n6753), .A2(n6752), .A3(n6751), .A4(n6750), .ZN(n6772) );
  AOI22D0 U2831 ( .A1(n6680), .A2(\mem[159][1] ), .B1(n6982), .B2(
        \mem[130][1] ), .ZN(n6758) );
  AOI22D0 U2832 ( .A1(n6888), .A2(\mem[128][1] ), .B1(n6891), .B2(
        \mem[154][1] ), .ZN(n6757) );
  AOI22D0 U2833 ( .A1(n6971), .A2(\mem[166][1] ), .B1(n6992), .B2(
        \mem[182][1] ), .ZN(n6756) );
  AOI22D0 U2834 ( .A1(n6926), .A2(\mem[129][1] ), .B1(n6754), .B2(
        \mem[133][1] ), .ZN(n6755) );
  ND4D0 U2835 ( .A1(n6758), .A2(n6757), .A3(n6756), .A4(n6755), .ZN(n6771) );
  AOI22D0 U2836 ( .A1(n6759), .A2(\mem[142][1] ), .B1(n6905), .B2(
        \mem[187][1] ), .ZN(n6764) );
  AOI22D0 U2837 ( .A1(n6927), .A2(\mem[153][1] ), .B1(n6760), .B2(
        \mem[173][1] ), .ZN(n6763) );
  AOI22D0 U2838 ( .A1(n6933), .A2(\mem[161][1] ), .B1(n6988), .B2(
        \mem[191][1] ), .ZN(n6761) );
  ND4D0 U2839 ( .A1(n6764), .A2(n6763), .A3(n6762), .A4(n6761), .ZN(n6770) );
  AOI22D0 U2840 ( .A1(n6952), .A2(\mem[150][1] ), .B1(n6958), .B2(
        \mem[145][1] ), .ZN(n6768) );
  AOI22D0 U2841 ( .A1(n6917), .A2(\mem[174][1] ), .B1(n6860), .B2(
        \mem[163][1] ), .ZN(n6767) );
  AOI22D0 U2842 ( .A1(n6863), .A2(\mem[183][1] ), .B1(n6990), .B2(
        \mem[140][1] ), .ZN(n6766) );
  AOI22D0 U2843 ( .A1(n6959), .A2(\mem[131][1] ), .B1(n6804), .B2(
        \mem[147][1] ), .ZN(n6765) );
  ND4D0 U2844 ( .A1(n6768), .A2(n6767), .A3(n6766), .A4(n6765), .ZN(n6769) );
  NR4D0 U2845 ( .A1(n6772), .A2(n6771), .A3(n6770), .A4(n6769), .ZN(n6801) );
  AOI22D0 U2846 ( .A1(n6773), .A2(\mem[164][1] ), .B1(n6964), .B2(
        \mem[158][1] ), .ZN(n6779) );
  AOI22D0 U2847 ( .A1(n6965), .A2(\mem[141][1] ), .B1(n6902), .B2(
        \mem[165][1] ), .ZN(n6778) );
  AOI22D0 U2848 ( .A1(n6957), .A2(\mem[185][1] ), .B1(n6912), .B2(
        \mem[184][1] ), .ZN(n6777) );
  AOI22D0 U2849 ( .A1(n6775), .A2(\mem[172][1] ), .B1(n6774), .B2(
        \mem[177][1] ), .ZN(n6776) );
  ND4D0 U2850 ( .A1(n6779), .A2(n6778), .A3(n6777), .A4(n6776), .ZN(n6799) );
  AOI22D0 U2851 ( .A1(n6880), .A2(\mem[139][1] ), .B1(n6954), .B2(
        \mem[138][1] ), .ZN(n6783) );
  AOI22D0 U2852 ( .A1(n6970), .A2(\mem[144][1] ), .B1(n6859), .B2(
        \mem[180][1] ), .ZN(n6782) );
  AOI22D0 U2853 ( .A1(n6819), .A2(\mem[189][1] ), .B1(n6922), .B2(
        \mem[157][1] ), .ZN(n6781) );
  AOI22D0 U2854 ( .A1(n6969), .A2(\mem[146][1] ), .B1(n6976), .B2(
        \mem[162][1] ), .ZN(n6780) );
  ND4D0 U2855 ( .A1(n6783), .A2(n6782), .A3(n6781), .A4(n6780), .ZN(n6798) );
  AOI22D0 U2856 ( .A1(n6989), .A2(\mem[134][1] ), .B1(n6883), .B2(
        \mem[176][1] ), .ZN(n6788) );
  AOI22D0 U2857 ( .A1(n6784), .A2(\mem[156][1] ), .B1(n6837), .B2(
        \mem[143][1] ), .ZN(n6786) );
  AOI22D0 U2858 ( .A1(n6870), .A2(\mem[188][1] ), .B1(n6862), .B2(
        \mem[168][1] ), .ZN(n6785) );
  ND4D0 U2859 ( .A1(n6788), .A2(n6787), .A3(n6786), .A4(n6785), .ZN(n6797) );
  AOI22D0 U2860 ( .A1(n6953), .A2(\mem[175][1] ), .B1(n6789), .B2(
        \mem[190][1] ), .ZN(n6795) );
  AOI22D0 U2861 ( .A1(n6802), .A2(\mem[152][1] ), .B1(n6790), .B2(
        \mem[155][1] ), .ZN(n6794) );
  AOI22D0 U2862 ( .A1(n6901), .A2(\mem[137][1] ), .B1(n6791), .B2(
        \mem[160][1] ), .ZN(n6793) );
  AOI22D0 U2863 ( .A1(n6967), .A2(\mem[167][1] ), .B1(n6966), .B2(
        \mem[178][1] ), .ZN(n6792) );
  ND4D0 U2864 ( .A1(n6795), .A2(n6794), .A3(n6793), .A4(n6792), .ZN(n6796) );
  NR4D0 U2865 ( .A1(n6799), .A2(n6798), .A3(n6797), .A4(n6796), .ZN(n6800) );
  CKND2D0 U2866 ( .A1(n6801), .A2(n6800), .ZN(n6950) );
  AOI22D0 U2867 ( .A1(n6802), .A2(\mem[24][1] ), .B1(n6916), .B2(\mem[21][1] ), 
        .ZN(n6808) );
  AOI22D0 U2868 ( .A1(n6803), .A2(\mem[55][1] ), .B1(n6966), .B2(\mem[50][1] ), 
        .ZN(n6807) );
  AOI22D0 U2869 ( .A1(n6905), .A2(\mem[59][1] ), .B1(n6804), .B2(\mem[19][1] ), 
        .ZN(n6806) );
  AOI22D0 U2870 ( .A1(n6913), .A2(\mem[27][1] ), .B1(n6903), .B2(\mem[51][1] ), 
        .ZN(n6805) );
  ND4D0 U2871 ( .A1(n6808), .A2(n6807), .A3(n6806), .A4(n6805), .ZN(n6827) );
  AOI22D0 U2872 ( .A1(n6879), .A2(\mem[58][1] ), .B1(n6995), .B2(\mem[23][1] ), 
        .ZN(n6813) );
  AOI22D0 U2873 ( .A1(n6953), .A2(\mem[47][1] ), .B1(n6892), .B2(\mem[44][1] ), 
        .ZN(n6812) );
  AOI22D0 U2874 ( .A1(n6809), .A2(\mem[9][1] ), .B1(n6935), .B2(\mem[63][1] ), 
        .ZN(n6811) );
  AOI22D0 U2875 ( .A1(n6889), .A2(\mem[28][1] ), .B1(n6982), .B2(\mem[2][1] ), 
        .ZN(n6810) );
  ND4D0 U2876 ( .A1(n6813), .A2(n6812), .A3(n6811), .A4(n6810), .ZN(n6826) );
  AOI22D0 U2877 ( .A1(n6952), .A2(\mem[22][1] ), .B1(n6923), .B2(\mem[34][1] ), 
        .ZN(n6817) );
  AOI22D0 U2878 ( .A1(n6880), .A2(\mem[11][1] ), .B1(n6814), .B2(\mem[1][1] ), 
        .ZN(n6816) );
  AOI22D0 U2879 ( .A1(n6969), .A2(\mem[18][1] ), .B1(n6906), .B2(\mem[12][1] ), 
        .ZN(n6815) );
  ND4D0 U2880 ( .A1(n6818), .A2(n6817), .A3(n6816), .A4(n6815), .ZN(n6825) );
  AOI22D0 U2881 ( .A1(n6819), .A2(\mem[61][1] ), .B1(n6977), .B2(\mem[33][1] ), 
        .ZN(n6823) );
  AOI22D0 U2882 ( .A1(n6883), .A2(\mem[48][1] ), .B1(n6956), .B2(\mem[40][1] ), 
        .ZN(n6822) );
  AOI22D0 U2883 ( .A1(n6860), .A2(\mem[35][1] ), .B1(n6869), .B2(\mem[49][1] ), 
        .ZN(n6821) );
  AOI22D0 U2884 ( .A1(n6868), .A2(\mem[43][1] ), .B1(n6881), .B2(\mem[16][1] ), 
        .ZN(n6820) );
  ND4D0 U2885 ( .A1(n6823), .A2(n6822), .A3(n6821), .A4(n6820), .ZN(n6824) );
  NR4D0 U2886 ( .A1(n6827), .A2(n6826), .A3(n6825), .A4(n6824), .ZN(n6858) );
  AOI22D0 U2887 ( .A1(n6873), .A2(\mem[30][1] ), .B1(n6828), .B2(\mem[56][1] ), 
        .ZN(n6834) );
  AOI22D0 U2888 ( .A1(n6830), .A2(\mem[7][1] ), .B1(n6829), .B2(\mem[38][1] ), 
        .ZN(n6833) );
  AOI22D0 U2889 ( .A1(n6917), .A2(\mem[46][1] ), .B1(n6871), .B2(\mem[57][1] ), 
        .ZN(n6832) );
  AOI22D0 U2890 ( .A1(n6994), .A2(\mem[62][1] ), .B1(n6968), .B2(\mem[41][1] ), 
        .ZN(n6831) );
  ND4D0 U2891 ( .A1(n6834), .A2(n6833), .A3(n6832), .A4(n6831), .ZN(n6855) );
  AOI22D0 U2892 ( .A1(n6981), .A2(\mem[60][1] ), .B1(n6835), .B2(\mem[4][1] ), 
        .ZN(n6841) );
  AOI22D0 U2893 ( .A1(n6872), .A2(\mem[6][1] ), .B1(n6936), .B2(\mem[17][1] ), 
        .ZN(n6840) );
  AOI22D0 U2894 ( .A1(n6890), .A2(\mem[36][1] ), .B1(n6836), .B2(\mem[10][1] ), 
        .ZN(n6839) );
  AOI22D0 U2895 ( .A1(n6991), .A2(\mem[20][1] ), .B1(n6888), .B2(\mem[0][1] ), 
        .ZN(n6846) );
  AOI22D0 U2896 ( .A1(n6925), .A2(\mem[45][1] ), .B1(n6978), .B2(\mem[8][1] ), 
        .ZN(n6845) );
  AOI22D0 U2897 ( .A1(n6993), .A2(\mem[53][1] ), .B1(n6859), .B2(\mem[52][1] ), 
        .ZN(n6844) );
  AOI22D0 U2898 ( .A1(n6842), .A2(\mem[26][1] ), .B1(n6992), .B2(\mem[54][1] ), 
        .ZN(n6843) );
  ND4D0 U2899 ( .A1(n6846), .A2(n6845), .A3(n6844), .A4(n6843), .ZN(n6853) );
  AOI22D0 U2900 ( .A1(n6907), .A2(\mem[3][1] ), .B1(n6979), .B2(\mem[14][1] ), 
        .ZN(n6851) );
  AOI22D0 U2901 ( .A1(n6680), .A2(\mem[31][1] ), .B1(n6902), .B2(\mem[37][1] ), 
        .ZN(n6850) );
  AOI22D0 U2902 ( .A1(n6847), .A2(\mem[25][1] ), .B1(n6924), .B2(\mem[32][1] ), 
        .ZN(n6849) );
  AOI22D0 U2903 ( .A1(n6874), .A2(\mem[42][1] ), .B1(n6965), .B2(\mem[13][1] ), 
        .ZN(n6848) );
  ND4D0 U2904 ( .A1(n6851), .A2(n6850), .A3(n6849), .A4(n6848), .ZN(n6852) );
  NR4D0 U2905 ( .A1(n6855), .A2(n6854), .A3(n6853), .A4(n6852), .ZN(n6857) );
  AOI21D0 U2906 ( .A1(n6858), .A2(n6857), .B(n6856), .ZN(n6949) );
  AOI22D0 U2907 ( .A1(n6860), .A2(\mem[227][1] ), .B1(n6859), .B2(
        \mem[244][1] ), .ZN(n6867) );
  AOI22D0 U2908 ( .A1(n6969), .A2(\mem[210][1] ), .B1(n6978), .B2(
        \mem[200][1] ), .ZN(n6866) );
  AOI22D0 U2909 ( .A1(n6861), .A2(\mem[196][1] ), .B1(n6992), .B2(
        \mem[246][1] ), .ZN(n6865) );
  AOI22D0 U2910 ( .A1(n6863), .A2(\mem[247][1] ), .B1(n6862), .B2(
        \mem[232][1] ), .ZN(n6864) );
  ND4D0 U2911 ( .A1(n6867), .A2(n6866), .A3(n6865), .A4(n6864), .ZN(n6900) );
  AOI22D0 U2912 ( .A1(n6868), .A2(\mem[235][1] ), .B1(n6968), .B2(
        \mem[233][1] ), .ZN(n6878) );
  AOI22D0 U2913 ( .A1(n6870), .A2(\mem[252][1] ), .B1(n6869), .B2(
        \mem[241][1] ), .ZN(n6877) );
  AOI22D0 U2914 ( .A1(n6874), .A2(\mem[234][1] ), .B1(n6873), .B2(
        \mem[222][1] ), .ZN(n6875) );
  ND4D0 U2915 ( .A1(n6878), .A2(n6877), .A3(n6876), .A4(n6875), .ZN(n6899) );
  AOI22D0 U2916 ( .A1(n6953), .A2(\mem[239][1] ), .B1(n6879), .B2(
        \mem[250][1] ), .ZN(n6887) );
  AOI22D0 U2917 ( .A1(n6880), .A2(\mem[203][1] ), .B1(n6994), .B2(
        \mem[254][1] ), .ZN(n6886) );
  AOI22D0 U2918 ( .A1(n6980), .A2(\mem[253][1] ), .B1(n6881), .B2(
        \mem[208][1] ), .ZN(n6885) );
  AOI22D0 U2919 ( .A1(n6883), .A2(\mem[240][1] ), .B1(n6882), .B2(
        \mem[207][1] ), .ZN(n6884) );
  ND4D0 U2920 ( .A1(n6887), .A2(n6886), .A3(n6885), .A4(n6884), .ZN(n6898) );
  AOI22D0 U2921 ( .A1(n6889), .A2(\mem[220][1] ), .B1(n6888), .B2(
        \mem[192][1] ), .ZN(n6896) );
  AOI22D0 U2922 ( .A1(n6680), .A2(\mem[223][1] ), .B1(n6995), .B2(
        \mem[215][1] ), .ZN(n6895) );
  AOI22D0 U2923 ( .A1(n6890), .A2(\mem[228][1] ), .B1(n6991), .B2(
        \mem[212][1] ), .ZN(n6894) );
  AOI22D0 U2924 ( .A1(n6892), .A2(\mem[236][1] ), .B1(n6891), .B2(
        \mem[218][1] ), .ZN(n6893) );
  ND4D0 U2925 ( .A1(n6896), .A2(n6895), .A3(n6894), .A4(n6893), .ZN(n6897) );
  NR4D0 U2926 ( .A1(n6900), .A2(n6899), .A3(n6898), .A4(n6897), .ZN(n6947) );
  AOI22D0 U2927 ( .A1(n6971), .A2(\mem[230][1] ), .B1(n6901), .B2(
        \mem[201][1] ), .ZN(n6911) );
  AOI22D0 U2928 ( .A1(n6903), .A2(\mem[243][1] ), .B1(n6902), .B2(
        \mem[229][1] ), .ZN(n6910) );
  AOI22D0 U2929 ( .A1(n6905), .A2(\mem[251][1] ), .B1(n6904), .B2(
        \mem[211][1] ), .ZN(n6909) );
  AOI22D0 U2930 ( .A1(n6907), .A2(\mem[195][1] ), .B1(n6906), .B2(
        \mem[204][1] ), .ZN(n6908) );
  ND4D0 U2931 ( .A1(n6911), .A2(n6910), .A3(n6909), .A4(n6908), .ZN(n6944) );
  AOI22D0 U2932 ( .A1(n6913), .A2(\mem[219][1] ), .B1(n6912), .B2(
        \mem[248][1] ), .ZN(n6921) );
  AOI22D0 U2933 ( .A1(n6979), .A2(\mem[206][1] ), .B1(n6915), .B2(
        \mem[205][1] ), .ZN(n6919) );
  AOI22D0 U2934 ( .A1(n6917), .A2(\mem[238][1] ), .B1(n6916), .B2(
        \mem[213][1] ), .ZN(n6918) );
  ND4D0 U2935 ( .A1(n6921), .A2(n6920), .A3(n6919), .A4(n6918), .ZN(n6943) );
  AOI22D0 U2936 ( .A1(n6923), .A2(\mem[226][1] ), .B1(n6922), .B2(
        \mem[221][1] ), .ZN(n6932) );
  AOI22D0 U2937 ( .A1(n6924), .A2(\mem[224][1] ), .B1(n6966), .B2(
        \mem[242][1] ), .ZN(n6931) );
  AOI22D0 U2938 ( .A1(n6926), .A2(\mem[193][1] ), .B1(n6925), .B2(
        \mem[237][1] ), .ZN(n6930) );
  AOI22D0 U2939 ( .A1(n6928), .A2(\mem[199][1] ), .B1(n6927), .B2(
        \mem[217][1] ), .ZN(n6929) );
  ND4D0 U2940 ( .A1(n6932), .A2(n6931), .A3(n6930), .A4(n6929), .ZN(n6942) );
  AOI22D0 U2941 ( .A1(n6952), .A2(\mem[214][1] ), .B1(n6933), .B2(
        \mem[225][1] ), .ZN(n6940) );
  AOI22D0 U2942 ( .A1(n6934), .A2(\mem[216][1] ), .B1(n6967), .B2(
        \mem[231][1] ), .ZN(n6939) );
  AOI22D0 U2943 ( .A1(n6954), .A2(\mem[202][1] ), .B1(n6935), .B2(
        \mem[255][1] ), .ZN(n6938) );
  AOI22D0 U2944 ( .A1(n6993), .A2(\mem[245][1] ), .B1(n6936), .B2(
        \mem[209][1] ), .ZN(n6937) );
  ND4D0 U2945 ( .A1(n6940), .A2(n6939), .A3(n6938), .A4(n6937), .ZN(n6941) );
  NR4D0 U2946 ( .A1(n6944), .A2(n6943), .A3(n6942), .A4(n6941), .ZN(n6946) );
  AOI21D0 U2947 ( .A1(n6947), .A2(n6946), .B(n6945), .ZN(n6948) );
  AOI211D0 U2948 ( .A1(n6951), .A2(n6950), .B(n6949), .C(n6948), .ZN(n7006) );
  AOI22D0 U2949 ( .A1(n6953), .A2(\mem[111][1] ), .B1(n6952), .B2(\mem[86][1] ), .ZN(n6963) );
  AOI22D0 U2950 ( .A1(n6955), .A2(\mem[85][1] ), .B1(n6954), .B2(\mem[74][1] ), 
        .ZN(n6962) );
  AOI22D0 U2951 ( .A1(n6957), .A2(\mem[121][1] ), .B1(n6956), .B2(
        \mem[104][1] ), .ZN(n6961) );
  AOI22D0 U2952 ( .A1(n6959), .A2(\mem[67][1] ), .B1(n6958), .B2(\mem[81][1] ), 
        .ZN(n6960) );
  ND4D0 U2953 ( .A1(n6963), .A2(n6962), .A3(n6961), .A4(n6960), .ZN(n7003) );
  AOI22D0 U2954 ( .A1(n6965), .A2(\mem[77][1] ), .B1(n6964), .B2(\mem[94][1] ), 
        .ZN(n6975) );
  AOI22D0 U2955 ( .A1(n6967), .A2(\mem[103][1] ), .B1(n6966), .B2(
        \mem[114][1] ), .ZN(n6974) );
  AOI22D0 U2956 ( .A1(n6971), .A2(\mem[102][1] ), .B1(n6970), .B2(\mem[80][1] ), .ZN(n6972) );
  ND4D0 U2957 ( .A1(n6975), .A2(n6974), .A3(n6973), .A4(n6972), .ZN(n7002) );
  AOI22D0 U2958 ( .A1(n6977), .A2(\mem[97][1] ), .B1(n6976), .B2(\mem[98][1] ), 
        .ZN(n6987) );
  AOI22D0 U2959 ( .A1(n6979), .A2(\mem[78][1] ), .B1(n6978), .B2(\mem[72][1] ), 
        .ZN(n6986) );
  AOI22D0 U2960 ( .A1(n6981), .A2(\mem[124][1] ), .B1(n6980), .B2(
        \mem[125][1] ), .ZN(n6985) );
  AOI22D0 U2961 ( .A1(n6983), .A2(\mem[112][1] ), .B1(n6982), .B2(\mem[66][1] ), .ZN(n6984) );
  AOI22D0 U2962 ( .A1(n6989), .A2(\mem[70][1] ), .B1(n6988), .B2(\mem[127][1] ), .ZN(n6999) );
  AOI22D0 U2963 ( .A1(n6991), .A2(\mem[84][1] ), .B1(n6990), .B2(\mem[76][1] ), 
        .ZN(n6998) );
  AOI22D0 U2964 ( .A1(n6993), .A2(\mem[117][1] ), .B1(n6992), .B2(
        \mem[118][1] ), .ZN(n6997) );
  AOI22D0 U2965 ( .A1(n6995), .A2(\mem[87][1] ), .B1(n6994), .B2(\mem[126][1] ), .ZN(n6996) );
  ND4D0 U2966 ( .A1(n6999), .A2(n6998), .A3(n6997), .A4(n6996), .ZN(n7000) );
  NR4D0 U2967 ( .A1(n7003), .A2(n7002), .A3(n7001), .A4(n7000), .ZN(n7005) );
  AOI32D0 U2968 ( .A1(n7007), .A2(n7006), .A3(n7005), .B1(n7004), .B2(n7006), 
        .ZN(dout[1]) );
  NR2D0 U2969 ( .A1(prog_addr[2]), .A2(prog_addr[1]), .ZN(n7032) );
  NR2D0 U2970 ( .A1(prog_addr[3]), .A2(prog_addr[0]), .ZN(n7022) );
  CKND2D0 U2971 ( .A1(n7032), .A2(n7022), .ZN(n7528) );
  INVD0 U2972 ( .I(prog_addr[5]), .ZN(n7187) );
  CKND2D0 U2973 ( .A1(prog_we), .A2(n7187), .ZN(n7458) );
  INVD0 U2974 ( .I(prog_addr[7]), .ZN(n7322) );
  CKND2D0 U2975 ( .A1(prog_we), .A2(n7322), .ZN(n7053) );
  NR2D0 U2976 ( .A1(prog_addr[4]), .A2(n7053), .ZN(n7221) );
  CKND2D0 U2977 ( .A1(n7324), .A2(n7221), .ZN(n7050) );
  INVD0 U2978 ( .I(n7008), .ZN(n7009) );
  OA22D0 U2979 ( .A1(n7009), .A2(prog_data[15]), .B1(\mem[0][15] ), .B2(n7008), 
        .Z(n4668) );
  OA22D0 U2980 ( .A1(n7009), .A2(prog_data[14]), .B1(\mem[0][14] ), .B2(n7008), 
        .Z(n4667) );
  OA22D0 U2981 ( .A1(n7009), .A2(prog_data[13]), .B1(\mem[0][13] ), .B2(n7008), 
        .Z(n4666) );
  OA22D0 U2982 ( .A1(n7009), .A2(prog_data[12]), .B1(\mem[0][12] ), .B2(n7008), 
        .Z(n4665) );
  OA22D0 U2983 ( .A1(n7009), .A2(prog_data[11]), .B1(\mem[0][11] ), .B2(n7008), 
        .Z(n4664) );
  OA22D0 U2984 ( .A1(n7009), .A2(prog_data[10]), .B1(\mem[0][10] ), .B2(n7008), 
        .Z(n4663) );
  OA22D0 U2985 ( .A1(n7009), .A2(prog_data[9]), .B1(\mem[0][9] ), .B2(n7008), 
        .Z(n4662) );
  OA22D0 U2986 ( .A1(n7009), .A2(prog_data[8]), .B1(\mem[0][8] ), .B2(n7008), 
        .Z(n4661) );
  OA22D0 U2987 ( .A1(n7009), .A2(prog_data[7]), .B1(\mem[0][7] ), .B2(n7008), 
        .Z(n4660) );
  OA22D0 U2988 ( .A1(n7009), .A2(prog_data[6]), .B1(\mem[0][6] ), .B2(n7008), 
        .Z(n4659) );
  OA22D0 U2989 ( .A1(n7009), .A2(prog_data[5]), .B1(\mem[0][5] ), .B2(n7008), 
        .Z(n4658) );
  OA22D0 U2990 ( .A1(n7009), .A2(prog_data[4]), .B1(\mem[0][4] ), .B2(n7008), 
        .Z(n4657) );
  OA22D0 U2991 ( .A1(n7009), .A2(prog_data[3]), .B1(\mem[0][3] ), .B2(n7008), 
        .Z(n4656) );
  OA22D0 U2992 ( .A1(n7009), .A2(prog_data[2]), .B1(\mem[0][2] ), .B2(n7008), 
        .Z(n4655) );
  OA22D0 U2993 ( .A1(n7009), .A2(prog_data[1]), .B1(\mem[0][1] ), .B2(n7008), 
        .Z(n4654) );
  OA22D0 U2994 ( .A1(n7009), .A2(prog_data[0]), .B1(\mem[0][0] ), .B2(n7008), 
        .Z(n4653) );
  INVD0 U2995 ( .I(prog_addr[0]), .ZN(n7030) );
  NR2D0 U2996 ( .A1(prog_addr[3]), .A2(n7030), .ZN(n7025) );
  CKND2D0 U2997 ( .A1(n7032), .A2(n7025), .ZN(n7531) );
  INVD0 U2998 ( .I(n7010), .ZN(n7011) );
  OA22D0 U2999 ( .A1(n7011), .A2(prog_data[15]), .B1(\mem[1][15] ), .B2(n7010), 
        .Z(n4652) );
  OA22D0 U3000 ( .A1(n7011), .A2(prog_data[14]), .B1(\mem[1][14] ), .B2(n7010), 
        .Z(n4651) );
  OA22D0 U3001 ( .A1(n7011), .A2(prog_data[13]), .B1(\mem[1][13] ), .B2(n7010), 
        .Z(n4650) );
  OA22D0 U3002 ( .A1(n7011), .A2(prog_data[12]), .B1(\mem[1][12] ), .B2(n7010), 
        .Z(n4649) );
  OA22D0 U3003 ( .A1(n7011), .A2(prog_data[11]), .B1(\mem[1][11] ), .B2(n7010), 
        .Z(n4648) );
  OA22D0 U3004 ( .A1(n7011), .A2(prog_data[10]), .B1(\mem[1][10] ), .B2(n7010), 
        .Z(n4647) );
  OA22D0 U3005 ( .A1(n7011), .A2(prog_data[9]), .B1(\mem[1][9] ), .B2(n7010), 
        .Z(n4646) );
  OA22D0 U3006 ( .A1(n7011), .A2(prog_data[8]), .B1(\mem[1][8] ), .B2(n7010), 
        .Z(n4645) );
  OA22D0 U3007 ( .A1(n7011), .A2(prog_data[7]), .B1(\mem[1][7] ), .B2(n7010), 
        .Z(n4644) );
  OA22D0 U3008 ( .A1(n7011), .A2(prog_data[6]), .B1(\mem[1][6] ), .B2(n7010), 
        .Z(n4643) );
  OA22D0 U3009 ( .A1(n7011), .A2(prog_data[5]), .B1(\mem[1][5] ), .B2(n7010), 
        .Z(n4642) );
  OA22D0 U3010 ( .A1(n7011), .A2(prog_data[4]), .B1(\mem[1][4] ), .B2(n7010), 
        .Z(n4641) );
  OA22D0 U3011 ( .A1(n7011), .A2(prog_data[3]), .B1(\mem[1][3] ), .B2(n7010), 
        .Z(n4640) );
  OA22D0 U3012 ( .A1(n7011), .A2(prog_data[2]), .B1(\mem[1][2] ), .B2(n7010), 
        .Z(n4639) );
  OA22D0 U3013 ( .A1(n7011), .A2(prog_data[1]), .B1(\mem[1][1] ), .B2(n7010), 
        .Z(n4638) );
  OA22D0 U3014 ( .A1(n7011), .A2(prog_data[0]), .B1(\mem[1][0] ), .B2(n7010), 
        .Z(n4637) );
  NR2D0 U3015 ( .A1(prog_addr[2]), .A2(n7020), .ZN(n7037) );
  CKND2D0 U3016 ( .A1(n7022), .A2(n7037), .ZN(n7534) );
  NR2D0 U3017 ( .A1(n7050), .A2(n7534), .ZN(n7012) );
  INVD0 U3018 ( .I(n7012), .ZN(n7013) );
  OA22D0 U3019 ( .A1(n7013), .A2(prog_data[15]), .B1(\mem[2][15] ), .B2(n7012), 
        .Z(n4636) );
  OA22D0 U3020 ( .A1(n7013), .A2(prog_data[14]), .B1(\mem[2][14] ), .B2(n7012), 
        .Z(n4635) );
  OA22D0 U3021 ( .A1(n7013), .A2(prog_data[13]), .B1(\mem[2][13] ), .B2(n7012), 
        .Z(n4634) );
  OA22D0 U3022 ( .A1(n7013), .A2(prog_data[12]), .B1(\mem[2][12] ), .B2(n7012), 
        .Z(n4633) );
  OA22D0 U3023 ( .A1(n7013), .A2(prog_data[11]), .B1(\mem[2][11] ), .B2(n7012), 
        .Z(n4632) );
  OA22D0 U3024 ( .A1(n7013), .A2(prog_data[10]), .B1(\mem[2][10] ), .B2(n7012), 
        .Z(n4631) );
  OA22D0 U3025 ( .A1(n7013), .A2(prog_data[9]), .B1(\mem[2][9] ), .B2(n7012), 
        .Z(n4630) );
  OA22D0 U3026 ( .A1(n7013), .A2(prog_data[8]), .B1(\mem[2][8] ), .B2(n7012), 
        .Z(n4629) );
  OA22D0 U3027 ( .A1(n7013), .A2(prog_data[7]), .B1(\mem[2][7] ), .B2(n7012), 
        .Z(n4628) );
  OA22D0 U3028 ( .A1(n7013), .A2(prog_data[6]), .B1(\mem[2][6] ), .B2(n7012), 
        .Z(n4627) );
  OA22D0 U3029 ( .A1(n7013), .A2(prog_data[5]), .B1(\mem[2][5] ), .B2(n7012), 
        .Z(n4626) );
  OA22D0 U3030 ( .A1(n7013), .A2(prog_data[4]), .B1(\mem[2][4] ), .B2(n7012), 
        .Z(n4625) );
  OA22D0 U3031 ( .A1(n7013), .A2(prog_data[3]), .B1(\mem[2][3] ), .B2(n7012), 
        .Z(n4624) );
  OA22D0 U3032 ( .A1(n7013), .A2(prog_data[2]), .B1(\mem[2][2] ), .B2(n7012), 
        .Z(n4623) );
  OA22D0 U3033 ( .A1(n7013), .A2(prog_data[1]), .B1(\mem[2][1] ), .B2(n7012), 
        .Z(n4622) );
  OA22D0 U3034 ( .A1(n7013), .A2(prog_data[0]), .B1(\mem[2][0] ), .B2(n7012), 
        .Z(n4621) );
  NR2D0 U3035 ( .A1(n7050), .A2(n7537), .ZN(n7014) );
  INVD0 U3036 ( .I(n7014), .ZN(n7015) );
  OA22D0 U3037 ( .A1(n7015), .A2(prog_data[15]), .B1(\mem[3][15] ), .B2(n7014), 
        .Z(n4620) );
  OA22D0 U3038 ( .A1(n7015), .A2(prog_data[14]), .B1(\mem[3][14] ), .B2(n7014), 
        .Z(n4619) );
  OA22D0 U3039 ( .A1(n7015), .A2(prog_data[13]), .B1(\mem[3][13] ), .B2(n7014), 
        .Z(n4618) );
  OA22D0 U3040 ( .A1(n7015), .A2(prog_data[12]), .B1(\mem[3][12] ), .B2(n7014), 
        .Z(n4617) );
  OA22D0 U3041 ( .A1(n7015), .A2(prog_data[11]), .B1(\mem[3][11] ), .B2(n7014), 
        .Z(n4616) );
  OA22D0 U3042 ( .A1(n7015), .A2(prog_data[10]), .B1(\mem[3][10] ), .B2(n7014), 
        .Z(n4615) );
  OA22D0 U3043 ( .A1(n7015), .A2(prog_data[9]), .B1(\mem[3][9] ), .B2(n7014), 
        .Z(n4614) );
  OA22D0 U3044 ( .A1(n7015), .A2(prog_data[8]), .B1(\mem[3][8] ), .B2(n7014), 
        .Z(n4613) );
  OA22D0 U3045 ( .A1(n7015), .A2(prog_data[7]), .B1(\mem[3][7] ), .B2(n7014), 
        .Z(n4612) );
  OA22D0 U3046 ( .A1(n7015), .A2(prog_data[6]), .B1(\mem[3][6] ), .B2(n7014), 
        .Z(n4611) );
  OA22D0 U3047 ( .A1(n7015), .A2(prog_data[5]), .B1(\mem[3][5] ), .B2(n7014), 
        .Z(n4610) );
  OA22D0 U3048 ( .A1(n7015), .A2(prog_data[4]), .B1(\mem[3][4] ), .B2(n7014), 
        .Z(n4609) );
  OA22D0 U3049 ( .A1(n7015), .A2(prog_data[3]), .B1(\mem[3][3] ), .B2(n7014), 
        .Z(n4608) );
  OA22D0 U3050 ( .A1(n7015), .A2(prog_data[2]), .B1(\mem[3][2] ), .B2(n7014), 
        .Z(n4607) );
  OA22D0 U3051 ( .A1(n7015), .A2(prog_data[1]), .B1(\mem[3][1] ), .B2(n7014), 
        .Z(n4606) );
  OA22D0 U3052 ( .A1(n7015), .A2(prog_data[0]), .B1(\mem[3][0] ), .B2(n7014), 
        .Z(n4605) );
  INVD0 U3053 ( .I(prog_addr[2]), .ZN(n7021) );
  NR2D0 U3054 ( .A1(prog_addr[1]), .A2(n7021), .ZN(n7042) );
  CKND2D0 U3055 ( .A1(n7022), .A2(n7042), .ZN(n7540) );
  NR2D0 U3056 ( .A1(n7050), .A2(n7540), .ZN(n7016) );
  INVD0 U3057 ( .I(n7016), .ZN(n7017) );
  OA22D0 U3058 ( .A1(n7017), .A2(prog_data[15]), .B1(\mem[4][15] ), .B2(n7016), 
        .Z(n4604) );
  OA22D0 U3059 ( .A1(n7017), .A2(prog_data[14]), .B1(\mem[4][14] ), .B2(n7016), 
        .Z(n4603) );
  OA22D0 U3060 ( .A1(n7017), .A2(prog_data[13]), .B1(\mem[4][13] ), .B2(n7016), 
        .Z(n4602) );
  OA22D0 U3061 ( .A1(n7017), .A2(prog_data[12]), .B1(\mem[4][12] ), .B2(n7016), 
        .Z(n4601) );
  OA22D0 U3062 ( .A1(n7017), .A2(prog_data[11]), .B1(\mem[4][11] ), .B2(n7016), 
        .Z(n4600) );
  OA22D0 U3063 ( .A1(n7017), .A2(prog_data[10]), .B1(\mem[4][10] ), .B2(n7016), 
        .Z(n4599) );
  OA22D0 U3064 ( .A1(n7017), .A2(prog_data[9]), .B1(\mem[4][9] ), .B2(n7016), 
        .Z(n4598) );
  OA22D0 U3065 ( .A1(n7017), .A2(prog_data[8]), .B1(\mem[4][8] ), .B2(n7016), 
        .Z(n4597) );
  OA22D0 U3066 ( .A1(n7017), .A2(prog_data[7]), .B1(\mem[4][7] ), .B2(n7016), 
        .Z(n4596) );
  OA22D0 U3067 ( .A1(n7017), .A2(prog_data[6]), .B1(\mem[4][6] ), .B2(n7016), 
        .Z(n4595) );
  OA22D0 U3068 ( .A1(n7017), .A2(prog_data[5]), .B1(\mem[4][5] ), .B2(n7016), 
        .Z(n4594) );
  OA22D0 U3069 ( .A1(n7017), .A2(prog_data[4]), .B1(\mem[4][4] ), .B2(n7016), 
        .Z(n4593) );
  OA22D0 U3070 ( .A1(n7017), .A2(prog_data[3]), .B1(\mem[4][3] ), .B2(n7016), 
        .Z(n4592) );
  OA22D0 U3071 ( .A1(n7017), .A2(prog_data[2]), .B1(\mem[4][2] ), .B2(n7016), 
        .Z(n4591) );
  OA22D0 U3072 ( .A1(n7017), .A2(prog_data[1]), .B1(\mem[4][1] ), .B2(n7016), 
        .Z(n4590) );
  OA22D0 U3073 ( .A1(n7017), .A2(prog_data[0]), .B1(\mem[4][0] ), .B2(n7016), 
        .Z(n4589) );
  CKND2D0 U3074 ( .A1(n7025), .A2(n7042), .ZN(n7543) );
  NR2D0 U3075 ( .A1(n7050), .A2(n7543), .ZN(n7018) );
  INVD0 U3076 ( .I(n7018), .ZN(n7019) );
  OA22D0 U3077 ( .A1(n7019), .A2(prog_data[15]), .B1(\mem[5][15] ), .B2(n7018), 
        .Z(n4588) );
  OA22D0 U3078 ( .A1(n7019), .A2(prog_data[14]), .B1(\mem[5][14] ), .B2(n7018), 
        .Z(n4587) );
  OA22D0 U3079 ( .A1(n7019), .A2(prog_data[13]), .B1(\mem[5][13] ), .B2(n7018), 
        .Z(n4586) );
  OA22D0 U3080 ( .A1(n7019), .A2(prog_data[12]), .B1(\mem[5][12] ), .B2(n7018), 
        .Z(n4585) );
  OA22D0 U3081 ( .A1(n7019), .A2(prog_data[11]), .B1(\mem[5][11] ), .B2(n7018), 
        .Z(n4584) );
  OA22D0 U3082 ( .A1(n7019), .A2(prog_data[10]), .B1(\mem[5][10] ), .B2(n7018), 
        .Z(n4583) );
  OA22D0 U3083 ( .A1(n7019), .A2(prog_data[9]), .B1(\mem[5][9] ), .B2(n7018), 
        .Z(n4582) );
  OA22D0 U3084 ( .A1(n7019), .A2(prog_data[8]), .B1(\mem[5][8] ), .B2(n7018), 
        .Z(n4581) );
  OA22D0 U3085 ( .A1(n7019), .A2(prog_data[7]), .B1(\mem[5][7] ), .B2(n7018), 
        .Z(n4580) );
  OA22D0 U3086 ( .A1(n7019), .A2(prog_data[6]), .B1(\mem[5][6] ), .B2(n7018), 
        .Z(n4579) );
  OA22D0 U3087 ( .A1(n7019), .A2(prog_data[5]), .B1(\mem[5][5] ), .B2(n7018), 
        .Z(n4578) );
  OA22D0 U3088 ( .A1(n7019), .A2(prog_data[4]), .B1(\mem[5][4] ), .B2(n7018), 
        .Z(n4577) );
  OA22D0 U3089 ( .A1(n7019), .A2(prog_data[3]), .B1(\mem[5][3] ), .B2(n7018), 
        .Z(n4576) );
  OA22D0 U3090 ( .A1(n7019), .A2(prog_data[2]), .B1(\mem[5][2] ), .B2(n7018), 
        .Z(n4575) );
  OA22D0 U3091 ( .A1(n7019), .A2(prog_data[1]), .B1(\mem[5][1] ), .B2(n7018), 
        .Z(n4574) );
  OA22D0 U3092 ( .A1(n7019), .A2(prog_data[0]), .B1(\mem[5][0] ), .B2(n7018), 
        .Z(n4573) );
  NR2D0 U3093 ( .A1(n7021), .A2(n7020), .ZN(n7049) );
  CKND2D0 U3094 ( .A1(n7022), .A2(n7049), .ZN(n7546) );
  NR2D0 U3095 ( .A1(n7050), .A2(n7546), .ZN(n7023) );
  INVD0 U3096 ( .I(n7023), .ZN(n7024) );
  OA22D0 U3097 ( .A1(n7024), .A2(prog_data[15]), .B1(\mem[6][15] ), .B2(n7023), 
        .Z(n4572) );
  OA22D0 U3098 ( .A1(n7024), .A2(prog_data[14]), .B1(\mem[6][14] ), .B2(n7023), 
        .Z(n4571) );
  OA22D0 U3099 ( .A1(n7024), .A2(prog_data[13]), .B1(\mem[6][13] ), .B2(n7023), 
        .Z(n4570) );
  OA22D0 U3100 ( .A1(n7024), .A2(prog_data[12]), .B1(\mem[6][12] ), .B2(n7023), 
        .Z(n4569) );
  OA22D0 U3101 ( .A1(n7024), .A2(prog_data[11]), .B1(\mem[6][11] ), .B2(n7023), 
        .Z(n4568) );
  OA22D0 U3102 ( .A1(n7024), .A2(prog_data[10]), .B1(\mem[6][10] ), .B2(n7023), 
        .Z(n4567) );
  OA22D0 U3103 ( .A1(n7024), .A2(prog_data[9]), .B1(\mem[6][9] ), .B2(n7023), 
        .Z(n4566) );
  OA22D0 U3104 ( .A1(n7024), .A2(prog_data[8]), .B1(\mem[6][8] ), .B2(n7023), 
        .Z(n4565) );
  OA22D0 U3105 ( .A1(n7024), .A2(prog_data[7]), .B1(\mem[6][7] ), .B2(n7023), 
        .Z(n4564) );
  OA22D0 U3106 ( .A1(n7024), .A2(prog_data[6]), .B1(\mem[6][6] ), .B2(n7023), 
        .Z(n4563) );
  OA22D0 U3107 ( .A1(n7024), .A2(prog_data[5]), .B1(\mem[6][5] ), .B2(n7023), 
        .Z(n4562) );
  OA22D0 U3108 ( .A1(n7024), .A2(prog_data[4]), .B1(\mem[6][4] ), .B2(n7023), 
        .Z(n4561) );
  OA22D0 U3109 ( .A1(n7024), .A2(prog_data[3]), .B1(\mem[6][3] ), .B2(n7023), 
        .Z(n4560) );
  OA22D0 U3110 ( .A1(n7024), .A2(prog_data[2]), .B1(\mem[6][2] ), .B2(n7023), 
        .Z(n4559) );
  OA22D0 U3111 ( .A1(n7024), .A2(prog_data[1]), .B1(\mem[6][1] ), .B2(n7023), 
        .Z(n4558) );
  OA22D0 U3112 ( .A1(n7024), .A2(prog_data[0]), .B1(\mem[6][0] ), .B2(n7023), 
        .Z(n4557) );
  CKND2D0 U3113 ( .A1(n7025), .A2(n7049), .ZN(n7549) );
  NR2D0 U3114 ( .A1(n7050), .A2(n7549), .ZN(n7026) );
  INVD0 U3115 ( .I(n7026), .ZN(n7027) );
  OA22D0 U3116 ( .A1(n7027), .A2(prog_data[15]), .B1(\mem[7][15] ), .B2(n7026), 
        .Z(n4556) );
  OA22D0 U3117 ( .A1(n7027), .A2(prog_data[14]), .B1(\mem[7][14] ), .B2(n7026), 
        .Z(n4555) );
  OA22D0 U3118 ( .A1(n7027), .A2(prog_data[13]), .B1(\mem[7][13] ), .B2(n7026), 
        .Z(n4554) );
  OA22D0 U3119 ( .A1(n7027), .A2(prog_data[12]), .B1(\mem[7][12] ), .B2(n7026), 
        .Z(n4553) );
  OA22D0 U3120 ( .A1(n7027), .A2(prog_data[11]), .B1(\mem[7][11] ), .B2(n7026), 
        .Z(n4552) );
  OA22D0 U3121 ( .A1(n7027), .A2(prog_data[10]), .B1(\mem[7][10] ), .B2(n7026), 
        .Z(n4551) );
  OA22D0 U3122 ( .A1(n7027), .A2(prog_data[9]), .B1(\mem[7][9] ), .B2(n7026), 
        .Z(n4550) );
  OA22D0 U3123 ( .A1(n7027), .A2(prog_data[8]), .B1(\mem[7][8] ), .B2(n7026), 
        .Z(n4549) );
  OA22D0 U3124 ( .A1(n7027), .A2(prog_data[7]), .B1(\mem[7][7] ), .B2(n7026), 
        .Z(n4548) );
  OA22D0 U3125 ( .A1(n7027), .A2(prog_data[6]), .B1(\mem[7][6] ), .B2(n7026), 
        .Z(n4547) );
  OA22D0 U3126 ( .A1(n7027), .A2(prog_data[5]), .B1(\mem[7][5] ), .B2(n7026), 
        .Z(n4546) );
  OA22D0 U3127 ( .A1(n7027), .A2(prog_data[4]), .B1(\mem[7][4] ), .B2(n7026), 
        .Z(n4545) );
  OA22D0 U3128 ( .A1(n7027), .A2(prog_data[3]), .B1(\mem[7][3] ), .B2(n7026), 
        .Z(n4544) );
  OA22D0 U3129 ( .A1(n7027), .A2(prog_data[2]), .B1(\mem[7][2] ), .B2(n7026), 
        .Z(n4543) );
  OA22D0 U3130 ( .A1(n7027), .A2(prog_data[1]), .B1(\mem[7][1] ), .B2(n7026), 
        .Z(n4542) );
  OA22D0 U3131 ( .A1(n7027), .A2(prog_data[0]), .B1(\mem[7][0] ), .B2(n7026), 
        .Z(n4541) );
  INVD0 U3132 ( .I(prog_addr[3]), .ZN(n7031) );
  NR2D0 U3133 ( .A1(prog_addr[0]), .A2(n7031), .ZN(n7045) );
  CKND2D0 U3134 ( .A1(n7032), .A2(n7045), .ZN(n7552) );
  NR2D0 U3135 ( .A1(n7050), .A2(n7552), .ZN(n7028) );
  INVD0 U3136 ( .I(n7028), .ZN(n7029) );
  OA22D0 U3137 ( .A1(n7029), .A2(prog_data[15]), .B1(\mem[8][15] ), .B2(n7028), 
        .Z(n4540) );
  OA22D0 U3138 ( .A1(n7029), .A2(prog_data[14]), .B1(\mem[8][14] ), .B2(n7028), 
        .Z(n4539) );
  OA22D0 U3139 ( .A1(n7029), .A2(prog_data[13]), .B1(\mem[8][13] ), .B2(n7028), 
        .Z(n4538) );
  OA22D0 U3140 ( .A1(n7029), .A2(prog_data[12]), .B1(\mem[8][12] ), .B2(n7028), 
        .Z(n4537) );
  OA22D0 U3141 ( .A1(n7029), .A2(prog_data[11]), .B1(\mem[8][11] ), .B2(n7028), 
        .Z(n4536) );
  OA22D0 U3142 ( .A1(n7029), .A2(prog_data[10]), .B1(\mem[8][10] ), .B2(n7028), 
        .Z(n4535) );
  OA22D0 U3143 ( .A1(n7029), .A2(prog_data[9]), .B1(\mem[8][9] ), .B2(n7028), 
        .Z(n4534) );
  OA22D0 U3144 ( .A1(n7029), .A2(prog_data[8]), .B1(\mem[8][8] ), .B2(n7028), 
        .Z(n4533) );
  OA22D0 U3145 ( .A1(n7029), .A2(prog_data[7]), .B1(\mem[8][7] ), .B2(n7028), 
        .Z(n4532) );
  OA22D0 U3146 ( .A1(n7029), .A2(prog_data[6]), .B1(\mem[8][6] ), .B2(n7028), 
        .Z(n4531) );
  OA22D0 U3147 ( .A1(n7029), .A2(prog_data[5]), .B1(\mem[8][5] ), .B2(n7028), 
        .Z(n4530) );
  OA22D0 U3148 ( .A1(n7029), .A2(prog_data[4]), .B1(\mem[8][4] ), .B2(n7028), 
        .Z(n4529) );
  OA22D0 U3149 ( .A1(n7029), .A2(prog_data[3]), .B1(\mem[8][3] ), .B2(n7028), 
        .Z(n4528) );
  OA22D0 U3150 ( .A1(n7029), .A2(prog_data[2]), .B1(\mem[8][2] ), .B2(n7028), 
        .Z(n4527) );
  OA22D0 U3151 ( .A1(n7029), .A2(prog_data[1]), .B1(\mem[8][1] ), .B2(n7028), 
        .Z(n4526) );
  OA22D0 U3152 ( .A1(n7029), .A2(prog_data[0]), .B1(\mem[8][0] ), .B2(n7028), 
        .Z(n4525) );
  NR2D0 U3153 ( .A1(n7031), .A2(n7030), .ZN(n7048) );
  CKND2D0 U3154 ( .A1(n7032), .A2(n7048), .ZN(n7555) );
  NR2D0 U3155 ( .A1(n7050), .A2(n7555), .ZN(n7033) );
  OA22D0 U3156 ( .A1(n7034), .A2(prog_data[15]), .B1(\mem[9][15] ), .B2(n7033), 
        .Z(n4524) );
  OA22D0 U3157 ( .A1(n7034), .A2(prog_data[14]), .B1(\mem[9][14] ), .B2(n7033), 
        .Z(n4523) );
  OA22D0 U3158 ( .A1(n7034), .A2(prog_data[13]), .B1(\mem[9][13] ), .B2(n7033), 
        .Z(n4522) );
  OA22D0 U3159 ( .A1(n7034), .A2(prog_data[12]), .B1(\mem[9][12] ), .B2(n7033), 
        .Z(n4521) );
  OA22D0 U3160 ( .A1(n7034), .A2(prog_data[11]), .B1(\mem[9][11] ), .B2(n7033), 
        .Z(n4520) );
  OA22D0 U3161 ( .A1(n7034), .A2(prog_data[10]), .B1(\mem[9][10] ), .B2(n7033), 
        .Z(n4519) );
  OA22D0 U3162 ( .A1(n7034), .A2(prog_data[9]), .B1(\mem[9][9] ), .B2(n7033), 
        .Z(n4518) );
  OA22D0 U3163 ( .A1(n7034), .A2(prog_data[8]), .B1(\mem[9][8] ), .B2(n7033), 
        .Z(n4517) );
  OA22D0 U3164 ( .A1(n7034), .A2(prog_data[7]), .B1(\mem[9][7] ), .B2(n7033), 
        .Z(n4516) );
  OA22D0 U3165 ( .A1(n7034), .A2(prog_data[6]), .B1(\mem[9][6] ), .B2(n7033), 
        .Z(n4515) );
  OA22D0 U3166 ( .A1(n7034), .A2(prog_data[5]), .B1(\mem[9][5] ), .B2(n7033), 
        .Z(n4514) );
  OA22D0 U3167 ( .A1(n7034), .A2(prog_data[4]), .B1(\mem[9][4] ), .B2(n7033), 
        .Z(n4513) );
  OA22D0 U3168 ( .A1(n7034), .A2(prog_data[3]), .B1(\mem[9][3] ), .B2(n7033), 
        .Z(n4512) );
  OA22D0 U3169 ( .A1(n7034), .A2(prog_data[2]), .B1(\mem[9][2] ), .B2(n7033), 
        .Z(n4511) );
  OA22D0 U3170 ( .A1(n7034), .A2(prog_data[1]), .B1(\mem[9][1] ), .B2(n7033), 
        .Z(n4510) );
  OA22D0 U3171 ( .A1(n7034), .A2(prog_data[0]), .B1(\mem[9][0] ), .B2(n7033), 
        .Z(n4509) );
  CKND2D0 U3172 ( .A1(n7037), .A2(n7045), .ZN(n7558) );
  NR2D0 U3173 ( .A1(n7050), .A2(n7558), .ZN(n7035) );
  INVD0 U3174 ( .I(n7035), .ZN(n7036) );
  OA22D0 U3175 ( .A1(n7036), .A2(prog_data[15]), .B1(\mem[10][15] ), .B2(n7035), .Z(n4508) );
  OA22D0 U3176 ( .A1(n7036), .A2(prog_data[14]), .B1(\mem[10][14] ), .B2(n7035), .Z(n4507) );
  OA22D0 U3177 ( .A1(n7036), .A2(prog_data[13]), .B1(\mem[10][13] ), .B2(n7035), .Z(n4506) );
  OA22D0 U3178 ( .A1(n7036), .A2(prog_data[12]), .B1(\mem[10][12] ), .B2(n7035), .Z(n4505) );
  OA22D0 U3179 ( .A1(n7036), .A2(prog_data[11]), .B1(\mem[10][11] ), .B2(n7035), .Z(n4504) );
  OA22D0 U3180 ( .A1(n7036), .A2(prog_data[10]), .B1(\mem[10][10] ), .B2(n7035), .Z(n4503) );
  OA22D0 U3181 ( .A1(n7036), .A2(prog_data[9]), .B1(\mem[10][9] ), .B2(n7035), 
        .Z(n4502) );
  OA22D0 U3182 ( .A1(n7036), .A2(prog_data[8]), .B1(\mem[10][8] ), .B2(n7035), 
        .Z(n4501) );
  OA22D0 U3183 ( .A1(n7036), .A2(prog_data[7]), .B1(\mem[10][7] ), .B2(n7035), 
        .Z(n4500) );
  OA22D0 U3184 ( .A1(n7036), .A2(prog_data[6]), .B1(\mem[10][6] ), .B2(n7035), 
        .Z(n4499) );
  OA22D0 U3185 ( .A1(n7036), .A2(prog_data[5]), .B1(\mem[10][5] ), .B2(n7035), 
        .Z(n4498) );
  OA22D0 U3186 ( .A1(n7036), .A2(prog_data[4]), .B1(\mem[10][4] ), .B2(n7035), 
        .Z(n4497) );
  OA22D0 U3187 ( .A1(n7036), .A2(prog_data[3]), .B1(\mem[10][3] ), .B2(n7035), 
        .Z(n4496) );
  OA22D0 U3188 ( .A1(n7036), .A2(prog_data[2]), .B1(\mem[10][2] ), .B2(n7035), 
        .Z(n4495) );
  OA22D0 U3189 ( .A1(n7036), .A2(prog_data[1]), .B1(\mem[10][1] ), .B2(n7035), 
        .Z(n4494) );
  OA22D0 U3190 ( .A1(n7036), .A2(prog_data[0]), .B1(\mem[10][0] ), .B2(n7035), 
        .Z(n4493) );
  CKND2D0 U3191 ( .A1(n7037), .A2(n7048), .ZN(n7561) );
  NR2D0 U3192 ( .A1(n7050), .A2(n7561), .ZN(n7038) );
  INVD0 U3193 ( .I(n7038), .ZN(n7039) );
  OA22D0 U3194 ( .A1(n7039), .A2(prog_data[15]), .B1(\mem[11][15] ), .B2(n7038), .Z(n4492) );
  OA22D0 U3195 ( .A1(n7039), .A2(prog_data[14]), .B1(\mem[11][14] ), .B2(n7038), .Z(n4491) );
  OA22D0 U3196 ( .A1(n7039), .A2(prog_data[13]), .B1(\mem[11][13] ), .B2(n7038), .Z(n4490) );
  OA22D0 U3197 ( .A1(n7039), .A2(prog_data[12]), .B1(\mem[11][12] ), .B2(n7038), .Z(n4489) );
  OA22D0 U3198 ( .A1(n7039), .A2(prog_data[11]), .B1(\mem[11][11] ), .B2(n7038), .Z(n4488) );
  OA22D0 U3199 ( .A1(n7039), .A2(prog_data[10]), .B1(\mem[11][10] ), .B2(n7038), .Z(n4487) );
  OA22D0 U3200 ( .A1(n7039), .A2(prog_data[9]), .B1(\mem[11][9] ), .B2(n7038), 
        .Z(n4486) );
  OA22D0 U3201 ( .A1(n7039), .A2(prog_data[8]), .B1(\mem[11][8] ), .B2(n7038), 
        .Z(n4485) );
  OA22D0 U3202 ( .A1(n7039), .A2(prog_data[7]), .B1(\mem[11][7] ), .B2(n7038), 
        .Z(n4484) );
  OA22D0 U3203 ( .A1(n7039), .A2(prog_data[6]), .B1(\mem[11][6] ), .B2(n7038), 
        .Z(n4483) );
  OA22D0 U3204 ( .A1(n7039), .A2(prog_data[5]), .B1(\mem[11][5] ), .B2(n7038), 
        .Z(n4482) );
  OA22D0 U3205 ( .A1(n7039), .A2(prog_data[4]), .B1(\mem[11][4] ), .B2(n7038), 
        .Z(n4481) );
  OA22D0 U3206 ( .A1(n7039), .A2(prog_data[3]), .B1(\mem[11][3] ), .B2(n7038), 
        .Z(n4480) );
  OA22D0 U3207 ( .A1(n7039), .A2(prog_data[2]), .B1(\mem[11][2] ), .B2(n7038), 
        .Z(n4479) );
  OA22D0 U3208 ( .A1(n7039), .A2(prog_data[1]), .B1(\mem[11][1] ), .B2(n7038), 
        .Z(n4478) );
  OA22D0 U3209 ( .A1(n7039), .A2(prog_data[0]), .B1(\mem[11][0] ), .B2(n7038), 
        .Z(n4477) );
  CKND2D0 U3210 ( .A1(n7042), .A2(n7045), .ZN(n7564) );
  NR2D0 U3211 ( .A1(n7050), .A2(n7564), .ZN(n7040) );
  INVD0 U3212 ( .I(n7040), .ZN(n7041) );
  OA22D0 U3213 ( .A1(n7041), .A2(prog_data[15]), .B1(\mem[12][15] ), .B2(n7040), .Z(n4476) );
  OA22D0 U3214 ( .A1(n7041), .A2(prog_data[14]), .B1(\mem[12][14] ), .B2(n7040), .Z(n4475) );
  OA22D0 U3215 ( .A1(n7041), .A2(prog_data[13]), .B1(\mem[12][13] ), .B2(n7040), .Z(n4474) );
  OA22D0 U3216 ( .A1(n7041), .A2(prog_data[12]), .B1(\mem[12][12] ), .B2(n7040), .Z(n4473) );
  OA22D0 U3217 ( .A1(n7041), .A2(prog_data[11]), .B1(\mem[12][11] ), .B2(n7040), .Z(n4472) );
  OA22D0 U3218 ( .A1(n7041), .A2(prog_data[10]), .B1(\mem[12][10] ), .B2(n7040), .Z(n4471) );
  OA22D0 U3219 ( .A1(n7041), .A2(prog_data[9]), .B1(\mem[12][9] ), .B2(n7040), 
        .Z(n4470) );
  OA22D0 U3220 ( .A1(n7041), .A2(prog_data[8]), .B1(\mem[12][8] ), .B2(n7040), 
        .Z(n4469) );
  OA22D0 U3221 ( .A1(n7041), .A2(prog_data[7]), .B1(\mem[12][7] ), .B2(n7040), 
        .Z(n4468) );
  OA22D0 U3222 ( .A1(n7041), .A2(prog_data[6]), .B1(\mem[12][6] ), .B2(n7040), 
        .Z(n4467) );
  OA22D0 U3223 ( .A1(n7041), .A2(prog_data[5]), .B1(\mem[12][5] ), .B2(n7040), 
        .Z(n4466) );
  OA22D0 U3224 ( .A1(n7041), .A2(prog_data[4]), .B1(\mem[12][4] ), .B2(n7040), 
        .Z(n4465) );
  OA22D0 U3225 ( .A1(n7041), .A2(prog_data[3]), .B1(\mem[12][3] ), .B2(n7040), 
        .Z(n4464) );
  OA22D0 U3226 ( .A1(n7041), .A2(prog_data[2]), .B1(\mem[12][2] ), .B2(n7040), 
        .Z(n4463) );
  OA22D0 U3227 ( .A1(n7041), .A2(prog_data[1]), .B1(\mem[12][1] ), .B2(n7040), 
        .Z(n4462) );
  OA22D0 U3228 ( .A1(n7041), .A2(prog_data[0]), .B1(\mem[12][0] ), .B2(n7040), 
        .Z(n4461) );
  CKND2D0 U3229 ( .A1(n7042), .A2(n7048), .ZN(n7567) );
  NR2D0 U3230 ( .A1(n7050), .A2(n7567), .ZN(n7043) );
  INVD0 U3231 ( .I(n7043), .ZN(n7044) );
  OA22D0 U3232 ( .A1(n7044), .A2(prog_data[15]), .B1(\mem[13][15] ), .B2(n7043), .Z(n4460) );
  OA22D0 U3233 ( .A1(n7044), .A2(prog_data[14]), .B1(\mem[13][14] ), .B2(n7043), .Z(n4459) );
  OA22D0 U3234 ( .A1(n7044), .A2(prog_data[13]), .B1(\mem[13][13] ), .B2(n7043), .Z(n4458) );
  OA22D0 U3235 ( .A1(n7044), .A2(prog_data[12]), .B1(\mem[13][12] ), .B2(n7043), .Z(n4457) );
  OA22D0 U3236 ( .A1(n7044), .A2(prog_data[11]), .B1(\mem[13][11] ), .B2(n7043), .Z(n4456) );
  OA22D0 U3237 ( .A1(n7044), .A2(prog_data[10]), .B1(\mem[13][10] ), .B2(n7043), .Z(n4455) );
  OA22D0 U3238 ( .A1(n7044), .A2(prog_data[9]), .B1(\mem[13][9] ), .B2(n7043), 
        .Z(n4454) );
  OA22D0 U3239 ( .A1(n7044), .A2(prog_data[8]), .B1(\mem[13][8] ), .B2(n7043), 
        .Z(n4453) );
  OA22D0 U3240 ( .A1(n7044), .A2(prog_data[7]), .B1(\mem[13][7] ), .B2(n7043), 
        .Z(n4452) );
  OA22D0 U3241 ( .A1(n7044), .A2(prog_data[6]), .B1(\mem[13][6] ), .B2(n7043), 
        .Z(n4451) );
  OA22D0 U3242 ( .A1(n7044), .A2(prog_data[5]), .B1(\mem[13][5] ), .B2(n7043), 
        .Z(n4450) );
  OA22D0 U3243 ( .A1(n7044), .A2(prog_data[4]), .B1(\mem[13][4] ), .B2(n7043), 
        .Z(n4449) );
  OA22D0 U3244 ( .A1(n7044), .A2(prog_data[3]), .B1(\mem[13][3] ), .B2(n7043), 
        .Z(n4448) );
  OA22D0 U3245 ( .A1(n7044), .A2(prog_data[2]), .B1(\mem[13][2] ), .B2(n7043), 
        .Z(n4447) );
  OA22D0 U3246 ( .A1(n7044), .A2(prog_data[1]), .B1(\mem[13][1] ), .B2(n7043), 
        .Z(n4446) );
  OA22D0 U3247 ( .A1(n7044), .A2(prog_data[0]), .B1(\mem[13][0] ), .B2(n7043), 
        .Z(n4445) );
  CKND2D0 U3248 ( .A1(n7049), .A2(n7045), .ZN(n7570) );
  NR2D0 U3249 ( .A1(n7050), .A2(n7570), .ZN(n7046) );
  INVD0 U3250 ( .I(n7046), .ZN(n7047) );
  OA22D0 U3251 ( .A1(n7047), .A2(prog_data[15]), .B1(\mem[14][15] ), .B2(n7046), .Z(n4444) );
  OA22D0 U3252 ( .A1(n7047), .A2(prog_data[14]), .B1(\mem[14][14] ), .B2(n7046), .Z(n4443) );
  OA22D0 U3253 ( .A1(n7047), .A2(prog_data[13]), .B1(\mem[14][13] ), .B2(n7046), .Z(n4442) );
  OA22D0 U3254 ( .A1(n7047), .A2(prog_data[12]), .B1(\mem[14][12] ), .B2(n7046), .Z(n4441) );
  OA22D0 U3255 ( .A1(n7047), .A2(prog_data[11]), .B1(\mem[14][11] ), .B2(n7046), .Z(n4440) );
  OA22D0 U3256 ( .A1(n7047), .A2(prog_data[10]), .B1(\mem[14][10] ), .B2(n7046), .Z(n4439) );
  OA22D0 U3257 ( .A1(n7047), .A2(prog_data[9]), .B1(\mem[14][9] ), .B2(n7046), 
        .Z(n4438) );
  OA22D0 U3258 ( .A1(n7047), .A2(prog_data[8]), .B1(\mem[14][8] ), .B2(n7046), 
        .Z(n4437) );
  OA22D0 U3259 ( .A1(n7047), .A2(prog_data[7]), .B1(\mem[14][7] ), .B2(n7046), 
        .Z(n4436) );
  OA22D0 U3260 ( .A1(n7047), .A2(prog_data[6]), .B1(\mem[14][6] ), .B2(n7046), 
        .Z(n4435) );
  OA22D0 U3261 ( .A1(n7047), .A2(prog_data[5]), .B1(\mem[14][5] ), .B2(n7046), 
        .Z(n4434) );
  OA22D0 U3262 ( .A1(n7047), .A2(prog_data[4]), .B1(\mem[14][4] ), .B2(n7046), 
        .Z(n4433) );
  OA22D0 U3263 ( .A1(n7047), .A2(prog_data[3]), .B1(\mem[14][3] ), .B2(n7046), 
        .Z(n4432) );
  OA22D0 U3264 ( .A1(n7047), .A2(prog_data[2]), .B1(\mem[14][2] ), .B2(n7046), 
        .Z(n4431) );
  OA22D0 U3265 ( .A1(n7047), .A2(prog_data[1]), .B1(\mem[14][1] ), .B2(n7046), 
        .Z(n4430) );
  OA22D0 U3266 ( .A1(n7047), .A2(prog_data[0]), .B1(\mem[14][0] ), .B2(n7046), 
        .Z(n4429) );
  CKND2D0 U3267 ( .A1(n7049), .A2(n7048), .ZN(n7574) );
  NR2D0 U3268 ( .A1(n7050), .A2(n7574), .ZN(n7051) );
  INVD0 U3269 ( .I(n7051), .ZN(n7052) );
  OA22D0 U3270 ( .A1(n7052), .A2(prog_data[15]), .B1(\mem[15][15] ), .B2(n7051), .Z(n4428) );
  OA22D0 U3271 ( .A1(n7052), .A2(prog_data[14]), .B1(\mem[15][14] ), .B2(n7051), .Z(n4427) );
  OA22D0 U3272 ( .A1(n7052), .A2(prog_data[13]), .B1(\mem[15][13] ), .B2(n7051), .Z(n4426) );
  OA22D0 U3273 ( .A1(n7052), .A2(prog_data[12]), .B1(\mem[15][12] ), .B2(n7051), .Z(n4425) );
  OA22D0 U3274 ( .A1(n7052), .A2(prog_data[11]), .B1(\mem[15][11] ), .B2(n7051), .Z(n4424) );
  OA22D0 U3275 ( .A1(n7052), .A2(prog_data[10]), .B1(\mem[15][10] ), .B2(n7051), .Z(n4423) );
  OA22D0 U3276 ( .A1(n7052), .A2(prog_data[9]), .B1(\mem[15][9] ), .B2(n7051), 
        .Z(n4422) );
  OA22D0 U3277 ( .A1(n7052), .A2(prog_data[8]), .B1(\mem[15][8] ), .B2(n7051), 
        .Z(n4421) );
  OA22D0 U3278 ( .A1(n7052), .A2(prog_data[7]), .B1(\mem[15][7] ), .B2(n7051), 
        .Z(n4420) );
  OA22D0 U3279 ( .A1(n7052), .A2(prog_data[6]), .B1(\mem[15][6] ), .B2(n7051), 
        .Z(n4419) );
  OA22D0 U3280 ( .A1(n7052), .A2(prog_data[5]), .B1(\mem[15][5] ), .B2(n7051), 
        .Z(n4418) );
  OA22D0 U3281 ( .A1(n7052), .A2(prog_data[4]), .B1(\mem[15][4] ), .B2(n7051), 
        .Z(n4417) );
  OA22D0 U3282 ( .A1(n7052), .A2(prog_data[3]), .B1(\mem[15][3] ), .B2(n7051), 
        .Z(n4416) );
  OA22D0 U3283 ( .A1(n7052), .A2(prog_data[2]), .B1(\mem[15][2] ), .B2(n7051), 
        .Z(n4415) );
  OA22D0 U3284 ( .A1(n7052), .A2(prog_data[1]), .B1(\mem[15][1] ), .B2(n7051), 
        .Z(n4414) );
  OA22D0 U3285 ( .A1(n7052), .A2(prog_data[0]), .B1(\mem[15][0] ), .B2(n7051), 
        .Z(n4413) );
  INVD0 U3286 ( .I(prog_addr[4]), .ZN(n7323) );
  NR2D0 U3287 ( .A1(n7323), .A2(n7053), .ZN(n7255) );
  CKND2D0 U3288 ( .A1(n7324), .A2(n7255), .ZN(n7084) );
  INVD0 U3289 ( .I(n7054), .ZN(n7055) );
  OA22D0 U3290 ( .A1(n7055), .A2(prog_data[15]), .B1(\mem[16][15] ), .B2(n7054), .Z(n4412) );
  OA22D0 U3291 ( .A1(n7055), .A2(prog_data[14]), .B1(\mem[16][14] ), .B2(n7054), .Z(n4411) );
  OA22D0 U3292 ( .A1(n7055), .A2(prog_data[13]), .B1(\mem[16][13] ), .B2(n7054), .Z(n4410) );
  OA22D0 U3293 ( .A1(n7055), .A2(prog_data[12]), .B1(\mem[16][12] ), .B2(n7054), .Z(n4409) );
  OA22D0 U3294 ( .A1(n7055), .A2(prog_data[11]), .B1(\mem[16][11] ), .B2(n7054), .Z(n4408) );
  OA22D0 U3295 ( .A1(n7055), .A2(prog_data[10]), .B1(\mem[16][10] ), .B2(n7054), .Z(n4407) );
  OA22D0 U3296 ( .A1(n7055), .A2(prog_data[9]), .B1(\mem[16][9] ), .B2(n7054), 
        .Z(n4406) );
  OA22D0 U3297 ( .A1(n7055), .A2(prog_data[8]), .B1(\mem[16][8] ), .B2(n7054), 
        .Z(n4405) );
  OA22D0 U3298 ( .A1(n7055), .A2(prog_data[7]), .B1(\mem[16][7] ), .B2(n7054), 
        .Z(n4404) );
  OA22D0 U3299 ( .A1(n7055), .A2(prog_data[6]), .B1(\mem[16][6] ), .B2(n7054), 
        .Z(n4403) );
  OA22D0 U3300 ( .A1(n7055), .A2(prog_data[5]), .B1(\mem[16][5] ), .B2(n7054), 
        .Z(n4402) );
  OA22D0 U3301 ( .A1(n7055), .A2(prog_data[4]), .B1(\mem[16][4] ), .B2(n7054), 
        .Z(n4401) );
  OA22D0 U3302 ( .A1(n7055), .A2(prog_data[3]), .B1(\mem[16][3] ), .B2(n7054), 
        .Z(n4400) );
  OA22D0 U3303 ( .A1(n7055), .A2(prog_data[2]), .B1(\mem[16][2] ), .B2(n7054), 
        .Z(n4399) );
  OA22D0 U3304 ( .A1(n7055), .A2(prog_data[1]), .B1(\mem[16][1] ), .B2(n7054), 
        .Z(n4398) );
  OA22D0 U3305 ( .A1(n7055), .A2(prog_data[0]), .B1(\mem[16][0] ), .B2(n7054), 
        .Z(n4397) );
  NR2D0 U3306 ( .A1(n7531), .A2(n7084), .ZN(n7056) );
  INVD0 U3307 ( .I(n7056), .ZN(n7057) );
  OA22D0 U3308 ( .A1(n7057), .A2(prog_data[15]), .B1(\mem[17][15] ), .B2(n7056), .Z(n4396) );
  OA22D0 U3309 ( .A1(n7057), .A2(prog_data[14]), .B1(\mem[17][14] ), .B2(n7056), .Z(n4395) );
  OA22D0 U3310 ( .A1(n7057), .A2(prog_data[13]), .B1(\mem[17][13] ), .B2(n7056), .Z(n4394) );
  OA22D0 U3311 ( .A1(n7057), .A2(prog_data[12]), .B1(\mem[17][12] ), .B2(n7056), .Z(n4393) );
  OA22D0 U3312 ( .A1(n7057), .A2(prog_data[11]), .B1(\mem[17][11] ), .B2(n7056), .Z(n4392) );
  OA22D0 U3313 ( .A1(n7057), .A2(prog_data[10]), .B1(\mem[17][10] ), .B2(n7056), .Z(n4391) );
  OA22D0 U3314 ( .A1(n7057), .A2(prog_data[9]), .B1(\mem[17][9] ), .B2(n7056), 
        .Z(n4390) );
  OA22D0 U3315 ( .A1(n7057), .A2(prog_data[8]), .B1(\mem[17][8] ), .B2(n7056), 
        .Z(n4389) );
  OA22D0 U3316 ( .A1(n7057), .A2(prog_data[7]), .B1(\mem[17][7] ), .B2(n7056), 
        .Z(n4388) );
  OA22D0 U3317 ( .A1(n7057), .A2(prog_data[6]), .B1(\mem[17][6] ), .B2(n7056), 
        .Z(n4387) );
  OA22D0 U3318 ( .A1(n7057), .A2(prog_data[5]), .B1(\mem[17][5] ), .B2(n7056), 
        .Z(n4386) );
  OA22D0 U3319 ( .A1(n7057), .A2(prog_data[4]), .B1(\mem[17][4] ), .B2(n7056), 
        .Z(n4385) );
  OA22D0 U3320 ( .A1(n7057), .A2(prog_data[3]), .B1(\mem[17][3] ), .B2(n7056), 
        .Z(n4384) );
  OA22D0 U3321 ( .A1(n7057), .A2(prog_data[2]), .B1(\mem[17][2] ), .B2(n7056), 
        .Z(n4383) );
  OA22D0 U3322 ( .A1(n7057), .A2(prog_data[1]), .B1(\mem[17][1] ), .B2(n7056), 
        .Z(n4382) );
  OA22D0 U3323 ( .A1(n7057), .A2(prog_data[0]), .B1(\mem[17][0] ), .B2(n7056), 
        .Z(n4381) );
  NR2D0 U3324 ( .A1(n7534), .A2(n7084), .ZN(n7058) );
  INVD0 U3325 ( .I(n7058), .ZN(n7059) );
  OA22D0 U3326 ( .A1(n7059), .A2(prog_data[15]), .B1(\mem[18][15] ), .B2(n7058), .Z(n4380) );
  OA22D0 U3327 ( .A1(n7059), .A2(prog_data[14]), .B1(\mem[18][14] ), .B2(n7058), .Z(n4379) );
  OA22D0 U3328 ( .A1(n7059), .A2(prog_data[13]), .B1(\mem[18][13] ), .B2(n7058), .Z(n4378) );
  OA22D0 U3329 ( .A1(n7059), .A2(prog_data[12]), .B1(\mem[18][12] ), .B2(n7058), .Z(n4377) );
  OA22D0 U3330 ( .A1(n7059), .A2(prog_data[11]), .B1(\mem[18][11] ), .B2(n7058), .Z(n4376) );
  OA22D0 U3331 ( .A1(n7059), .A2(prog_data[10]), .B1(\mem[18][10] ), .B2(n7058), .Z(n4375) );
  OA22D0 U3332 ( .A1(n7059), .A2(prog_data[9]), .B1(\mem[18][9] ), .B2(n7058), 
        .Z(n4374) );
  OA22D0 U3333 ( .A1(n7059), .A2(prog_data[8]), .B1(\mem[18][8] ), .B2(n7058), 
        .Z(n4373) );
  OA22D0 U3334 ( .A1(n7059), .A2(prog_data[7]), .B1(\mem[18][7] ), .B2(n7058), 
        .Z(n4372) );
  OA22D0 U3335 ( .A1(n7059), .A2(prog_data[6]), .B1(\mem[18][6] ), .B2(n7058), 
        .Z(n4371) );
  OA22D0 U3336 ( .A1(n7059), .A2(prog_data[5]), .B1(\mem[18][5] ), .B2(n7058), 
        .Z(n4370) );
  OA22D0 U3337 ( .A1(n7059), .A2(prog_data[4]), .B1(\mem[18][4] ), .B2(n7058), 
        .Z(n4369) );
  OA22D0 U3338 ( .A1(n7059), .A2(prog_data[3]), .B1(\mem[18][3] ), .B2(n7058), 
        .Z(n4368) );
  OA22D0 U3339 ( .A1(n7059), .A2(prog_data[2]), .B1(\mem[18][2] ), .B2(n7058), 
        .Z(n4367) );
  OA22D0 U3340 ( .A1(n7059), .A2(prog_data[1]), .B1(\mem[18][1] ), .B2(n7058), 
        .Z(n4366) );
  OA22D0 U3341 ( .A1(n7059), .A2(prog_data[0]), .B1(\mem[18][0] ), .B2(n7058), 
        .Z(n4365) );
  NR2D0 U3342 ( .A1(n7537), .A2(n7084), .ZN(n7060) );
  INVD0 U3343 ( .I(n7060), .ZN(n7061) );
  OA22D0 U3344 ( .A1(n7061), .A2(prog_data[15]), .B1(\mem[19][15] ), .B2(n7060), .Z(n4364) );
  OA22D0 U3345 ( .A1(n7061), .A2(prog_data[14]), .B1(\mem[19][14] ), .B2(n7060), .Z(n4363) );
  OA22D0 U3346 ( .A1(n7061), .A2(prog_data[13]), .B1(\mem[19][13] ), .B2(n7060), .Z(n4362) );
  OA22D0 U3347 ( .A1(n7061), .A2(prog_data[12]), .B1(\mem[19][12] ), .B2(n7060), .Z(n4361) );
  OA22D0 U3348 ( .A1(n7061), .A2(prog_data[11]), .B1(\mem[19][11] ), .B2(n7060), .Z(n4360) );
  OA22D0 U3349 ( .A1(n7061), .A2(prog_data[10]), .B1(\mem[19][10] ), .B2(n7060), .Z(n4359) );
  OA22D0 U3350 ( .A1(n7061), .A2(prog_data[9]), .B1(\mem[19][9] ), .B2(n7060), 
        .Z(n4358) );
  OA22D0 U3351 ( .A1(n7061), .A2(prog_data[8]), .B1(\mem[19][8] ), .B2(n7060), 
        .Z(n4357) );
  OA22D0 U3352 ( .A1(n7061), .A2(prog_data[7]), .B1(\mem[19][7] ), .B2(n7060), 
        .Z(n4356) );
  OA22D0 U3353 ( .A1(n7061), .A2(prog_data[6]), .B1(\mem[19][6] ), .B2(n7060), 
        .Z(n4355) );
  OA22D0 U3354 ( .A1(n7061), .A2(prog_data[5]), .B1(\mem[19][5] ), .B2(n7060), 
        .Z(n4354) );
  OA22D0 U3355 ( .A1(n7061), .A2(prog_data[4]), .B1(\mem[19][4] ), .B2(n7060), 
        .Z(n4353) );
  OA22D0 U3356 ( .A1(n7061), .A2(prog_data[3]), .B1(\mem[19][3] ), .B2(n7060), 
        .Z(n4352) );
  OA22D0 U3357 ( .A1(n7061), .A2(prog_data[2]), .B1(\mem[19][2] ), .B2(n7060), 
        .Z(n4351) );
  OA22D0 U3358 ( .A1(n7061), .A2(prog_data[1]), .B1(\mem[19][1] ), .B2(n7060), 
        .Z(n4350) );
  OA22D0 U3359 ( .A1(n7061), .A2(prog_data[0]), .B1(\mem[19][0] ), .B2(n7060), 
        .Z(n4349) );
  NR2D0 U3360 ( .A1(n7540), .A2(n7084), .ZN(n7062) );
  INVD0 U3361 ( .I(n7062), .ZN(n7063) );
  OA22D0 U3362 ( .A1(n7063), .A2(prog_data[15]), .B1(\mem[20][15] ), .B2(n7062), .Z(n4348) );
  OA22D0 U3363 ( .A1(n7063), .A2(prog_data[14]), .B1(\mem[20][14] ), .B2(n7062), .Z(n4347) );
  OA22D0 U3364 ( .A1(n7063), .A2(prog_data[13]), .B1(\mem[20][13] ), .B2(n7062), .Z(n4346) );
  OA22D0 U3365 ( .A1(n7063), .A2(prog_data[12]), .B1(\mem[20][12] ), .B2(n7062), .Z(n4345) );
  OA22D0 U3366 ( .A1(n7063), .A2(prog_data[11]), .B1(\mem[20][11] ), .B2(n7062), .Z(n4344) );
  OA22D0 U3367 ( .A1(n7063), .A2(prog_data[10]), .B1(\mem[20][10] ), .B2(n7062), .Z(n4343) );
  OA22D0 U3368 ( .A1(n7063), .A2(prog_data[9]), .B1(\mem[20][9] ), .B2(n7062), 
        .Z(n4342) );
  OA22D0 U3369 ( .A1(n7063), .A2(prog_data[8]), .B1(\mem[20][8] ), .B2(n7062), 
        .Z(n4341) );
  OA22D0 U3370 ( .A1(n7063), .A2(prog_data[7]), .B1(\mem[20][7] ), .B2(n7062), 
        .Z(n4340) );
  OA22D0 U3371 ( .A1(n7063), .A2(prog_data[6]), .B1(\mem[20][6] ), .B2(n7062), 
        .Z(n4339) );
  OA22D0 U3372 ( .A1(n7063), .A2(prog_data[5]), .B1(\mem[20][5] ), .B2(n7062), 
        .Z(n4338) );
  OA22D0 U3373 ( .A1(n7063), .A2(prog_data[4]), .B1(\mem[20][4] ), .B2(n7062), 
        .Z(n4337) );
  OA22D0 U3374 ( .A1(n7063), .A2(prog_data[3]), .B1(\mem[20][3] ), .B2(n7062), 
        .Z(n4336) );
  OA22D0 U3375 ( .A1(n7063), .A2(prog_data[2]), .B1(\mem[20][2] ), .B2(n7062), 
        .Z(n4335) );
  OA22D0 U3376 ( .A1(n7063), .A2(prog_data[1]), .B1(\mem[20][1] ), .B2(n7062), 
        .Z(n4334) );
  OA22D0 U3377 ( .A1(n7063), .A2(prog_data[0]), .B1(\mem[20][0] ), .B2(n7062), 
        .Z(n4333) );
  NR2D0 U3378 ( .A1(n7543), .A2(n7084), .ZN(n7064) );
  INVD0 U3379 ( .I(n7064), .ZN(n7065) );
  OA22D0 U3380 ( .A1(n7065), .A2(prog_data[15]), .B1(\mem[21][15] ), .B2(n7064), .Z(n4332) );
  OA22D0 U3381 ( .A1(n7065), .A2(prog_data[14]), .B1(\mem[21][14] ), .B2(n7064), .Z(n4331) );
  OA22D0 U3382 ( .A1(n7065), .A2(prog_data[13]), .B1(\mem[21][13] ), .B2(n7064), .Z(n4330) );
  OA22D0 U3383 ( .A1(n7065), .A2(prog_data[12]), .B1(\mem[21][12] ), .B2(n7064), .Z(n4329) );
  OA22D0 U3384 ( .A1(n7065), .A2(prog_data[11]), .B1(\mem[21][11] ), .B2(n7064), .Z(n4328) );
  OA22D0 U3385 ( .A1(n7065), .A2(prog_data[10]), .B1(\mem[21][10] ), .B2(n7064), .Z(n4327) );
  OA22D0 U3386 ( .A1(n7065), .A2(prog_data[9]), .B1(\mem[21][9] ), .B2(n7064), 
        .Z(n4326) );
  OA22D0 U3387 ( .A1(n7065), .A2(prog_data[8]), .B1(\mem[21][8] ), .B2(n7064), 
        .Z(n4325) );
  OA22D0 U3388 ( .A1(n7065), .A2(prog_data[7]), .B1(\mem[21][7] ), .B2(n7064), 
        .Z(n4324) );
  OA22D0 U3389 ( .A1(n7065), .A2(prog_data[6]), .B1(\mem[21][6] ), .B2(n7064), 
        .Z(n4323) );
  OA22D0 U3390 ( .A1(n7065), .A2(prog_data[5]), .B1(\mem[21][5] ), .B2(n7064), 
        .Z(n4322) );
  OA22D0 U3391 ( .A1(n7065), .A2(prog_data[4]), .B1(\mem[21][4] ), .B2(n7064), 
        .Z(n4321) );
  OA22D0 U3392 ( .A1(n7065), .A2(prog_data[3]), .B1(\mem[21][3] ), .B2(n7064), 
        .Z(n4320) );
  OA22D0 U3393 ( .A1(n7065), .A2(prog_data[2]), .B1(\mem[21][2] ), .B2(n7064), 
        .Z(n4319) );
  OA22D0 U3394 ( .A1(n7065), .A2(prog_data[1]), .B1(\mem[21][1] ), .B2(n7064), 
        .Z(n4318) );
  OA22D0 U3395 ( .A1(n7065), .A2(prog_data[0]), .B1(\mem[21][0] ), .B2(n7064), 
        .Z(n4317) );
  NR2D0 U3396 ( .A1(n7546), .A2(n7084), .ZN(n7066) );
  INVD0 U3397 ( .I(n7066), .ZN(n7067) );
  OA22D0 U3398 ( .A1(n7067), .A2(prog_data[15]), .B1(\mem[22][15] ), .B2(n7066), .Z(n4316) );
  OA22D0 U3399 ( .A1(n7067), .A2(prog_data[14]), .B1(\mem[22][14] ), .B2(n7066), .Z(n4315) );
  OA22D0 U3400 ( .A1(n7067), .A2(prog_data[13]), .B1(\mem[22][13] ), .B2(n7066), .Z(n4314) );
  OA22D0 U3401 ( .A1(n7067), .A2(prog_data[12]), .B1(\mem[22][12] ), .B2(n7066), .Z(n4313) );
  OA22D0 U3402 ( .A1(n7067), .A2(prog_data[11]), .B1(\mem[22][11] ), .B2(n7066), .Z(n4312) );
  OA22D0 U3403 ( .A1(n7067), .A2(prog_data[10]), .B1(\mem[22][10] ), .B2(n7066), .Z(n4311) );
  OA22D0 U3404 ( .A1(n7067), .A2(prog_data[9]), .B1(\mem[22][9] ), .B2(n7066), 
        .Z(n4310) );
  OA22D0 U3405 ( .A1(n7067), .A2(prog_data[8]), .B1(\mem[22][8] ), .B2(n7066), 
        .Z(n4309) );
  OA22D0 U3406 ( .A1(n7067), .A2(prog_data[7]), .B1(\mem[22][7] ), .B2(n7066), 
        .Z(n4308) );
  OA22D0 U3407 ( .A1(n7067), .A2(prog_data[6]), .B1(\mem[22][6] ), .B2(n7066), 
        .Z(n4307) );
  OA22D0 U3408 ( .A1(n7067), .A2(prog_data[5]), .B1(\mem[22][5] ), .B2(n7066), 
        .Z(n4306) );
  OA22D0 U3409 ( .A1(n7067), .A2(prog_data[4]), .B1(\mem[22][4] ), .B2(n7066), 
        .Z(n4305) );
  OA22D0 U3410 ( .A1(n7067), .A2(prog_data[3]), .B1(\mem[22][3] ), .B2(n7066), 
        .Z(n4304) );
  OA22D0 U3411 ( .A1(n7067), .A2(prog_data[2]), .B1(\mem[22][2] ), .B2(n7066), 
        .Z(n4303) );
  OA22D0 U3412 ( .A1(n7067), .A2(prog_data[1]), .B1(\mem[22][1] ), .B2(n7066), 
        .Z(n4302) );
  OA22D0 U3413 ( .A1(n7067), .A2(prog_data[0]), .B1(\mem[22][0] ), .B2(n7066), 
        .Z(n4301) );
  NR2D0 U3414 ( .A1(n7549), .A2(n7084), .ZN(n7068) );
  INVD0 U3415 ( .I(n7068), .ZN(n7069) );
  OA22D0 U3416 ( .A1(n7069), .A2(prog_data[15]), .B1(\mem[23][15] ), .B2(n7068), .Z(n4300) );
  OA22D0 U3417 ( .A1(n7069), .A2(prog_data[14]), .B1(\mem[23][14] ), .B2(n7068), .Z(n4299) );
  OA22D0 U3418 ( .A1(n7069), .A2(prog_data[13]), .B1(\mem[23][13] ), .B2(n7068), .Z(n4298) );
  OA22D0 U3419 ( .A1(n7069), .A2(prog_data[12]), .B1(\mem[23][12] ), .B2(n7068), .Z(n4297) );
  OA22D0 U3420 ( .A1(n7069), .A2(prog_data[11]), .B1(\mem[23][11] ), .B2(n7068), .Z(n4296) );
  OA22D0 U3421 ( .A1(n7069), .A2(prog_data[10]), .B1(\mem[23][10] ), .B2(n7068), .Z(n4295) );
  OA22D0 U3422 ( .A1(n7069), .A2(prog_data[9]), .B1(\mem[23][9] ), .B2(n7068), 
        .Z(n4294) );
  OA22D0 U3423 ( .A1(n7069), .A2(prog_data[8]), .B1(\mem[23][8] ), .B2(n7068), 
        .Z(n4293) );
  OA22D0 U3424 ( .A1(n7069), .A2(prog_data[7]), .B1(\mem[23][7] ), .B2(n7068), 
        .Z(n4292) );
  OA22D0 U3425 ( .A1(n7069), .A2(prog_data[6]), .B1(\mem[23][6] ), .B2(n7068), 
        .Z(n4291) );
  OA22D0 U3426 ( .A1(n7069), .A2(prog_data[5]), .B1(\mem[23][5] ), .B2(n7068), 
        .Z(n4290) );
  OA22D0 U3427 ( .A1(n7069), .A2(prog_data[4]), .B1(\mem[23][4] ), .B2(n7068), 
        .Z(n4289) );
  OA22D0 U3428 ( .A1(n7069), .A2(prog_data[3]), .B1(\mem[23][3] ), .B2(n7068), 
        .Z(n4288) );
  OA22D0 U3429 ( .A1(n7069), .A2(prog_data[2]), .B1(\mem[23][2] ), .B2(n7068), 
        .Z(n4287) );
  OA22D0 U3430 ( .A1(n7069), .A2(prog_data[1]), .B1(\mem[23][1] ), .B2(n7068), 
        .Z(n4286) );
  OA22D0 U3431 ( .A1(n7069), .A2(prog_data[0]), .B1(\mem[23][0] ), .B2(n7068), 
        .Z(n4285) );
  NR2D0 U3432 ( .A1(n7552), .A2(n7084), .ZN(n7070) );
  OA22D0 U3433 ( .A1(n7071), .A2(prog_data[15]), .B1(\mem[24][15] ), .B2(n7070), .Z(n4284) );
  OA22D0 U3434 ( .A1(n7071), .A2(prog_data[14]), .B1(\mem[24][14] ), .B2(n7070), .Z(n4283) );
  OA22D0 U3435 ( .A1(n7071), .A2(prog_data[13]), .B1(\mem[24][13] ), .B2(n7070), .Z(n4282) );
  OA22D0 U3436 ( .A1(n7071), .A2(prog_data[12]), .B1(\mem[24][12] ), .B2(n7070), .Z(n4281) );
  OA22D0 U3437 ( .A1(n7071), .A2(prog_data[11]), .B1(\mem[24][11] ), .B2(n7070), .Z(n4280) );
  OA22D0 U3438 ( .A1(n7071), .A2(prog_data[10]), .B1(\mem[24][10] ), .B2(n7070), .Z(n4279) );
  OA22D0 U3439 ( .A1(n7071), .A2(prog_data[9]), .B1(\mem[24][9] ), .B2(n7070), 
        .Z(n4278) );
  OA22D0 U3440 ( .A1(n7071), .A2(prog_data[8]), .B1(\mem[24][8] ), .B2(n7070), 
        .Z(n4277) );
  OA22D0 U3441 ( .A1(n7071), .A2(prog_data[7]), .B1(\mem[24][7] ), .B2(n7070), 
        .Z(n4276) );
  OA22D0 U3442 ( .A1(n7071), .A2(prog_data[6]), .B1(\mem[24][6] ), .B2(n7070), 
        .Z(n4275) );
  OA22D0 U3443 ( .A1(n7071), .A2(prog_data[5]), .B1(\mem[24][5] ), .B2(n7070), 
        .Z(n4274) );
  OA22D0 U3444 ( .A1(n7071), .A2(prog_data[4]), .B1(\mem[24][4] ), .B2(n7070), 
        .Z(n4273) );
  OA22D0 U3445 ( .A1(n7071), .A2(prog_data[3]), .B1(\mem[24][3] ), .B2(n7070), 
        .Z(n4272) );
  OA22D0 U3446 ( .A1(n7071), .A2(prog_data[2]), .B1(\mem[24][2] ), .B2(n7070), 
        .Z(n4271) );
  OA22D0 U3447 ( .A1(n7071), .A2(prog_data[1]), .B1(\mem[24][1] ), .B2(n7070), 
        .Z(n4270) );
  OA22D0 U3448 ( .A1(n7071), .A2(prog_data[0]), .B1(\mem[24][0] ), .B2(n7070), 
        .Z(n4269) );
  NR2D0 U3449 ( .A1(n7555), .A2(n7084), .ZN(n7072) );
  INVD0 U3450 ( .I(n7072), .ZN(n7073) );
  OA22D0 U3451 ( .A1(n7073), .A2(prog_data[15]), .B1(\mem[25][15] ), .B2(n7072), .Z(n4268) );
  OA22D0 U3452 ( .A1(n7073), .A2(prog_data[14]), .B1(\mem[25][14] ), .B2(n7072), .Z(n4267) );
  OA22D0 U3453 ( .A1(n7073), .A2(prog_data[13]), .B1(\mem[25][13] ), .B2(n7072), .Z(n4266) );
  OA22D0 U3454 ( .A1(n7073), .A2(prog_data[12]), .B1(\mem[25][12] ), .B2(n7072), .Z(n4265) );
  OA22D0 U3455 ( .A1(n7073), .A2(prog_data[11]), .B1(\mem[25][11] ), .B2(n7072), .Z(n4264) );
  OA22D0 U3456 ( .A1(n7073), .A2(prog_data[10]), .B1(\mem[25][10] ), .B2(n7072), .Z(n4263) );
  OA22D0 U3457 ( .A1(n7073), .A2(prog_data[9]), .B1(\mem[25][9] ), .B2(n7072), 
        .Z(n4262) );
  OA22D0 U3458 ( .A1(n7073), .A2(prog_data[8]), .B1(\mem[25][8] ), .B2(n7072), 
        .Z(n4261) );
  OA22D0 U3459 ( .A1(n7073), .A2(prog_data[7]), .B1(\mem[25][7] ), .B2(n7072), 
        .Z(n4260) );
  OA22D0 U3460 ( .A1(n7073), .A2(prog_data[6]), .B1(\mem[25][6] ), .B2(n7072), 
        .Z(n4259) );
  OA22D0 U3461 ( .A1(n7073), .A2(prog_data[5]), .B1(\mem[25][5] ), .B2(n7072), 
        .Z(n4258) );
  OA22D0 U3462 ( .A1(n7073), .A2(prog_data[4]), .B1(\mem[25][4] ), .B2(n7072), 
        .Z(n4257) );
  OA22D0 U3463 ( .A1(n7073), .A2(prog_data[3]), .B1(\mem[25][3] ), .B2(n7072), 
        .Z(n4256) );
  OA22D0 U3464 ( .A1(n7073), .A2(prog_data[2]), .B1(\mem[25][2] ), .B2(n7072), 
        .Z(n4255) );
  OA22D0 U3465 ( .A1(n7073), .A2(prog_data[1]), .B1(\mem[25][1] ), .B2(n7072), 
        .Z(n4254) );
  OA22D0 U3466 ( .A1(n7073), .A2(prog_data[0]), .B1(\mem[25][0] ), .B2(n7072), 
        .Z(n4253) );
  NR2D0 U3467 ( .A1(n7558), .A2(n7084), .ZN(n7074) );
  INVD0 U3468 ( .I(n7074), .ZN(n7075) );
  OA22D0 U3469 ( .A1(n7075), .A2(prog_data[15]), .B1(\mem[26][15] ), .B2(n7074), .Z(n4252) );
  OA22D0 U3470 ( .A1(n7075), .A2(prog_data[14]), .B1(\mem[26][14] ), .B2(n7074), .Z(n4251) );
  OA22D0 U3471 ( .A1(n7075), .A2(prog_data[13]), .B1(\mem[26][13] ), .B2(n7074), .Z(n4250) );
  OA22D0 U3472 ( .A1(n7075), .A2(prog_data[12]), .B1(\mem[26][12] ), .B2(n7074), .Z(n4249) );
  OA22D0 U3473 ( .A1(n7075), .A2(prog_data[11]), .B1(\mem[26][11] ), .B2(n7074), .Z(n4248) );
  OA22D0 U3474 ( .A1(n7075), .A2(prog_data[10]), .B1(\mem[26][10] ), .B2(n7074), .Z(n4247) );
  OA22D0 U3475 ( .A1(n7075), .A2(prog_data[9]), .B1(\mem[26][9] ), .B2(n7074), 
        .Z(n4246) );
  OA22D0 U3476 ( .A1(n7075), .A2(prog_data[8]), .B1(\mem[26][8] ), .B2(n7074), 
        .Z(n4245) );
  OA22D0 U3477 ( .A1(n7075), .A2(prog_data[7]), .B1(\mem[26][7] ), .B2(n7074), 
        .Z(n4244) );
  OA22D0 U3478 ( .A1(n7075), .A2(prog_data[6]), .B1(\mem[26][6] ), .B2(n7074), 
        .Z(n4243) );
  OA22D0 U3479 ( .A1(n7075), .A2(prog_data[5]), .B1(\mem[26][5] ), .B2(n7074), 
        .Z(n4242) );
  OA22D0 U3480 ( .A1(n7075), .A2(prog_data[4]), .B1(\mem[26][4] ), .B2(n7074), 
        .Z(n4241) );
  OA22D0 U3481 ( .A1(n7075), .A2(prog_data[3]), .B1(\mem[26][3] ), .B2(n7074), 
        .Z(n4240) );
  OA22D0 U3482 ( .A1(n7075), .A2(prog_data[2]), .B1(\mem[26][2] ), .B2(n7074), 
        .Z(n4239) );
  OA22D0 U3483 ( .A1(n7075), .A2(prog_data[1]), .B1(\mem[26][1] ), .B2(n7074), 
        .Z(n4238) );
  OA22D0 U3484 ( .A1(n7075), .A2(prog_data[0]), .B1(\mem[26][0] ), .B2(n7074), 
        .Z(n4237) );
  NR2D0 U3485 ( .A1(n7561), .A2(n7084), .ZN(n7076) );
  INVD0 U3486 ( .I(n7076), .ZN(n7077) );
  OA22D0 U3487 ( .A1(n7077), .A2(prog_data[15]), .B1(\mem[27][15] ), .B2(n7076), .Z(n4236) );
  OA22D0 U3488 ( .A1(n7077), .A2(prog_data[14]), .B1(\mem[27][14] ), .B2(n7076), .Z(n4235) );
  OA22D0 U3489 ( .A1(n7077), .A2(prog_data[13]), .B1(\mem[27][13] ), .B2(n7076), .Z(n4234) );
  OA22D0 U3490 ( .A1(n7077), .A2(prog_data[12]), .B1(\mem[27][12] ), .B2(n7076), .Z(n4233) );
  OA22D0 U3491 ( .A1(n7077), .A2(prog_data[11]), .B1(\mem[27][11] ), .B2(n7076), .Z(n4232) );
  OA22D0 U3492 ( .A1(n7077), .A2(prog_data[10]), .B1(\mem[27][10] ), .B2(n7076), .Z(n4231) );
  OA22D0 U3493 ( .A1(n7077), .A2(prog_data[9]), .B1(\mem[27][9] ), .B2(n7076), 
        .Z(n4230) );
  OA22D0 U3494 ( .A1(n7077), .A2(prog_data[8]), .B1(\mem[27][8] ), .B2(n7076), 
        .Z(n4229) );
  OA22D0 U3495 ( .A1(n7077), .A2(prog_data[7]), .B1(\mem[27][7] ), .B2(n7076), 
        .Z(n4228) );
  OA22D0 U3496 ( .A1(n7077), .A2(prog_data[6]), .B1(\mem[27][6] ), .B2(n7076), 
        .Z(n4227) );
  OA22D0 U3497 ( .A1(n7077), .A2(prog_data[5]), .B1(\mem[27][5] ), .B2(n7076), 
        .Z(n4226) );
  OA22D0 U3498 ( .A1(n7077), .A2(prog_data[4]), .B1(\mem[27][4] ), .B2(n7076), 
        .Z(n4225) );
  OA22D0 U3499 ( .A1(n7077), .A2(prog_data[3]), .B1(\mem[27][3] ), .B2(n7076), 
        .Z(n4224) );
  OA22D0 U3500 ( .A1(n7077), .A2(prog_data[2]), .B1(\mem[27][2] ), .B2(n7076), 
        .Z(n4223) );
  OA22D0 U3501 ( .A1(n7077), .A2(prog_data[1]), .B1(\mem[27][1] ), .B2(n7076), 
        .Z(n4222) );
  OA22D0 U3502 ( .A1(n7077), .A2(prog_data[0]), .B1(\mem[27][0] ), .B2(n7076), 
        .Z(n4221) );
  NR2D0 U3503 ( .A1(n7564), .A2(n7084), .ZN(n7078) );
  INVD0 U3504 ( .I(n7078), .ZN(n7079) );
  OA22D0 U3505 ( .A1(n7079), .A2(prog_data[15]), .B1(\mem[28][15] ), .B2(n7078), .Z(n4220) );
  OA22D0 U3506 ( .A1(n7079), .A2(prog_data[14]), .B1(\mem[28][14] ), .B2(n7078), .Z(n4219) );
  OA22D0 U3507 ( .A1(n7079), .A2(prog_data[13]), .B1(\mem[28][13] ), .B2(n7078), .Z(n4218) );
  OA22D0 U3508 ( .A1(n7079), .A2(prog_data[12]), .B1(\mem[28][12] ), .B2(n7078), .Z(n4217) );
  OA22D0 U3509 ( .A1(n7079), .A2(prog_data[11]), .B1(\mem[28][11] ), .B2(n7078), .Z(n4216) );
  OA22D0 U3510 ( .A1(n7079), .A2(prog_data[10]), .B1(\mem[28][10] ), .B2(n7078), .Z(n4215) );
  OA22D0 U3511 ( .A1(n7079), .A2(prog_data[9]), .B1(\mem[28][9] ), .B2(n7078), 
        .Z(n4214) );
  OA22D0 U3512 ( .A1(n7079), .A2(prog_data[8]), .B1(\mem[28][8] ), .B2(n7078), 
        .Z(n4213) );
  OA22D0 U3513 ( .A1(n7079), .A2(prog_data[7]), .B1(\mem[28][7] ), .B2(n7078), 
        .Z(n4212) );
  OA22D0 U3514 ( .A1(n7079), .A2(prog_data[6]), .B1(\mem[28][6] ), .B2(n7078), 
        .Z(n4211) );
  OA22D0 U3515 ( .A1(n7079), .A2(prog_data[5]), .B1(\mem[28][5] ), .B2(n7078), 
        .Z(n4210) );
  OA22D0 U3516 ( .A1(n7079), .A2(prog_data[4]), .B1(\mem[28][4] ), .B2(n7078), 
        .Z(n4209) );
  OA22D0 U3517 ( .A1(n7079), .A2(prog_data[3]), .B1(\mem[28][3] ), .B2(n7078), 
        .Z(n4208) );
  OA22D0 U3518 ( .A1(n7079), .A2(prog_data[2]), .B1(\mem[28][2] ), .B2(n7078), 
        .Z(n4207) );
  OA22D0 U3519 ( .A1(n7079), .A2(prog_data[1]), .B1(\mem[28][1] ), .B2(n7078), 
        .Z(n4206) );
  OA22D0 U3520 ( .A1(n7079), .A2(prog_data[0]), .B1(\mem[28][0] ), .B2(n7078), 
        .Z(n4205) );
  NR2D0 U3521 ( .A1(n7567), .A2(n7084), .ZN(n7080) );
  INVD0 U3522 ( .I(n7080), .ZN(n7081) );
  OA22D0 U3523 ( .A1(n7081), .A2(prog_data[15]), .B1(\mem[29][15] ), .B2(n7080), .Z(n4204) );
  OA22D0 U3524 ( .A1(n7081), .A2(prog_data[14]), .B1(\mem[29][14] ), .B2(n7080), .Z(n4203) );
  OA22D0 U3525 ( .A1(n7081), .A2(prog_data[13]), .B1(\mem[29][13] ), .B2(n7080), .Z(n4202) );
  OA22D0 U3526 ( .A1(n7081), .A2(prog_data[12]), .B1(\mem[29][12] ), .B2(n7080), .Z(n4201) );
  OA22D0 U3527 ( .A1(n7081), .A2(prog_data[11]), .B1(\mem[29][11] ), .B2(n7080), .Z(n4200) );
  OA22D0 U3528 ( .A1(n7081), .A2(prog_data[10]), .B1(\mem[29][10] ), .B2(n7080), .Z(n4199) );
  OA22D0 U3529 ( .A1(n7081), .A2(prog_data[9]), .B1(\mem[29][9] ), .B2(n7080), 
        .Z(n4198) );
  OA22D0 U3530 ( .A1(n7081), .A2(prog_data[8]), .B1(\mem[29][8] ), .B2(n7080), 
        .Z(n4197) );
  OA22D0 U3531 ( .A1(n7081), .A2(prog_data[7]), .B1(\mem[29][7] ), .B2(n7080), 
        .Z(n4196) );
  OA22D0 U3532 ( .A1(n7081), .A2(prog_data[6]), .B1(\mem[29][6] ), .B2(n7080), 
        .Z(n4195) );
  OA22D0 U3533 ( .A1(n7081), .A2(prog_data[5]), .B1(\mem[29][5] ), .B2(n7080), 
        .Z(n4194) );
  OA22D0 U3534 ( .A1(n7081), .A2(prog_data[4]), .B1(\mem[29][4] ), .B2(n7080), 
        .Z(n4193) );
  OA22D0 U3535 ( .A1(n7081), .A2(prog_data[3]), .B1(\mem[29][3] ), .B2(n7080), 
        .Z(n4192) );
  OA22D0 U3536 ( .A1(n7081), .A2(prog_data[2]), .B1(\mem[29][2] ), .B2(n7080), 
        .Z(n4191) );
  OA22D0 U3537 ( .A1(n7081), .A2(prog_data[1]), .B1(\mem[29][1] ), .B2(n7080), 
        .Z(n4190) );
  OA22D0 U3538 ( .A1(n7081), .A2(prog_data[0]), .B1(\mem[29][0] ), .B2(n7080), 
        .Z(n4189) );
  NR2D0 U3539 ( .A1(n7570), .A2(n7084), .ZN(n7082) );
  INVD0 U3540 ( .I(n7082), .ZN(n7083) );
  OA22D0 U3541 ( .A1(n7083), .A2(prog_data[15]), .B1(\mem[30][15] ), .B2(n7082), .Z(n4188) );
  OA22D0 U3542 ( .A1(n7083), .A2(prog_data[14]), .B1(\mem[30][14] ), .B2(n7082), .Z(n4187) );
  OA22D0 U3543 ( .A1(n7083), .A2(prog_data[13]), .B1(\mem[30][13] ), .B2(n7082), .Z(n4186) );
  OA22D0 U3544 ( .A1(n7083), .A2(prog_data[12]), .B1(\mem[30][12] ), .B2(n7082), .Z(n4185) );
  OA22D0 U3545 ( .A1(n7083), .A2(prog_data[11]), .B1(\mem[30][11] ), .B2(n7082), .Z(n4184) );
  OA22D0 U3546 ( .A1(n7083), .A2(prog_data[10]), .B1(\mem[30][10] ), .B2(n7082), .Z(n4183) );
  OA22D0 U3547 ( .A1(n7083), .A2(prog_data[9]), .B1(\mem[30][9] ), .B2(n7082), 
        .Z(n4182) );
  OA22D0 U3548 ( .A1(n7083), .A2(prog_data[8]), .B1(\mem[30][8] ), .B2(n7082), 
        .Z(n4181) );
  OA22D0 U3549 ( .A1(n7083), .A2(prog_data[7]), .B1(\mem[30][7] ), .B2(n7082), 
        .Z(n4180) );
  OA22D0 U3550 ( .A1(n7083), .A2(prog_data[6]), .B1(\mem[30][6] ), .B2(n7082), 
        .Z(n4179) );
  OA22D0 U3551 ( .A1(n7083), .A2(prog_data[5]), .B1(\mem[30][5] ), .B2(n7082), 
        .Z(n4178) );
  OA22D0 U3552 ( .A1(n7083), .A2(prog_data[4]), .B1(\mem[30][4] ), .B2(n7082), 
        .Z(n4177) );
  OA22D0 U3553 ( .A1(n7083), .A2(prog_data[3]), .B1(\mem[30][3] ), .B2(n7082), 
        .Z(n4176) );
  OA22D0 U3554 ( .A1(n7083), .A2(prog_data[2]), .B1(\mem[30][2] ), .B2(n7082), 
        .Z(n4175) );
  OA22D0 U3555 ( .A1(n7083), .A2(prog_data[1]), .B1(\mem[30][1] ), .B2(n7082), 
        .Z(n4174) );
  OA22D0 U3556 ( .A1(n7083), .A2(prog_data[0]), .B1(\mem[30][0] ), .B2(n7082), 
        .Z(n4173) );
  INVD0 U3557 ( .I(n7085), .ZN(n7086) );
  OA22D0 U3558 ( .A1(n7086), .A2(prog_data[15]), .B1(\mem[31][15] ), .B2(n7085), .Z(n4172) );
  OA22D0 U3559 ( .A1(n7086), .A2(prog_data[14]), .B1(\mem[31][14] ), .B2(n7085), .Z(n4171) );
  OA22D0 U3560 ( .A1(n7086), .A2(prog_data[13]), .B1(\mem[31][13] ), .B2(n7085), .Z(n4170) );
  OA22D0 U3561 ( .A1(n7086), .A2(prog_data[12]), .B1(\mem[31][12] ), .B2(n7085), .Z(n4169) );
  OA22D0 U3562 ( .A1(n7086), .A2(prog_data[11]), .B1(\mem[31][11] ), .B2(n7085), .Z(n4168) );
  OA22D0 U3563 ( .A1(n7086), .A2(prog_data[10]), .B1(\mem[31][10] ), .B2(n7085), .Z(n4167) );
  OA22D0 U3564 ( .A1(n7086), .A2(prog_data[9]), .B1(\mem[31][9] ), .B2(n7085), 
        .Z(n4166) );
  OA22D0 U3565 ( .A1(n7086), .A2(prog_data[8]), .B1(\mem[31][8] ), .B2(n7085), 
        .Z(n4165) );
  OA22D0 U3566 ( .A1(n7086), .A2(prog_data[7]), .B1(\mem[31][7] ), .B2(n7085), 
        .Z(n4164) );
  OA22D0 U3567 ( .A1(n7086), .A2(prog_data[6]), .B1(\mem[31][6] ), .B2(n7085), 
        .Z(n4163) );
  OA22D0 U3568 ( .A1(n7086), .A2(prog_data[5]), .B1(\mem[31][5] ), .B2(n7085), 
        .Z(n4162) );
  OA22D0 U3569 ( .A1(n7086), .A2(prog_data[4]), .B1(\mem[31][4] ), .B2(n7085), 
        .Z(n4161) );
  OA22D0 U3570 ( .A1(n7086), .A2(prog_data[3]), .B1(\mem[31][3] ), .B2(n7085), 
        .Z(n4160) );
  OA22D0 U3571 ( .A1(n7086), .A2(prog_data[2]), .B1(\mem[31][2] ), .B2(n7085), 
        .Z(n4159) );
  OA22D0 U3572 ( .A1(n7086), .A2(prog_data[1]), .B1(\mem[31][1] ), .B2(n7085), 
        .Z(n4158) );
  OA22D0 U3573 ( .A1(n7086), .A2(prog_data[0]), .B1(\mem[31][0] ), .B2(n7085), 
        .Z(n4157) );
  NR2D0 U3574 ( .A1(prog_addr[6]), .A2(n7187), .ZN(n7120) );
  CKND2D0 U3575 ( .A1(n7221), .A2(n7120), .ZN(n7117) );
  NR2D0 U3576 ( .A1(n7528), .A2(n7117), .ZN(n7087) );
  INVD0 U3577 ( .I(n7087), .ZN(n7088) );
  OA22D0 U3578 ( .A1(n7088), .A2(prog_data[15]), .B1(\mem[32][15] ), .B2(n7087), .Z(n4156) );
  OA22D0 U3579 ( .A1(n7088), .A2(prog_data[14]), .B1(\mem[32][14] ), .B2(n7087), .Z(n4155) );
  OA22D0 U3580 ( .A1(n7088), .A2(prog_data[13]), .B1(\mem[32][13] ), .B2(n7087), .Z(n4154) );
  OA22D0 U3581 ( .A1(n7088), .A2(prog_data[12]), .B1(\mem[32][12] ), .B2(n7087), .Z(n4153) );
  OA22D0 U3582 ( .A1(n7088), .A2(prog_data[11]), .B1(\mem[32][11] ), .B2(n7087), .Z(n4152) );
  OA22D0 U3583 ( .A1(n7088), .A2(prog_data[10]), .B1(\mem[32][10] ), .B2(n7087), .Z(n4151) );
  OA22D0 U3584 ( .A1(n7088), .A2(prog_data[9]), .B1(\mem[32][9] ), .B2(n7087), 
        .Z(n4150) );
  OA22D0 U3585 ( .A1(n7088), .A2(prog_data[8]), .B1(\mem[32][8] ), .B2(n7087), 
        .Z(n4149) );
  OA22D0 U3586 ( .A1(n7088), .A2(prog_data[7]), .B1(\mem[32][7] ), .B2(n7087), 
        .Z(n4148) );
  OA22D0 U3587 ( .A1(n7088), .A2(prog_data[6]), .B1(\mem[32][6] ), .B2(n7087), 
        .Z(n4147) );
  OA22D0 U3588 ( .A1(n7088), .A2(prog_data[5]), .B1(\mem[32][5] ), .B2(n7087), 
        .Z(n4146) );
  OA22D0 U3589 ( .A1(n7088), .A2(prog_data[4]), .B1(\mem[32][4] ), .B2(n7087), 
        .Z(n4145) );
  OA22D0 U3590 ( .A1(n7088), .A2(prog_data[3]), .B1(\mem[32][3] ), .B2(n7087), 
        .Z(n4144) );
  OA22D0 U3591 ( .A1(n7088), .A2(prog_data[2]), .B1(\mem[32][2] ), .B2(n7087), 
        .Z(n4143) );
  OA22D0 U3592 ( .A1(n7088), .A2(prog_data[1]), .B1(\mem[32][1] ), .B2(n7087), 
        .Z(n4142) );
  OA22D0 U3593 ( .A1(n7088), .A2(prog_data[0]), .B1(\mem[32][0] ), .B2(n7087), 
        .Z(n4141) );
  NR2D0 U3594 ( .A1(n7531), .A2(n7117), .ZN(n7089) );
  INVD0 U3595 ( .I(n7089), .ZN(n7090) );
  OA22D0 U3596 ( .A1(n7090), .A2(prog_data[15]), .B1(\mem[33][15] ), .B2(n7089), .Z(n4140) );
  OA22D0 U3597 ( .A1(n7090), .A2(prog_data[14]), .B1(\mem[33][14] ), .B2(n7089), .Z(n4139) );
  OA22D0 U3598 ( .A1(n7090), .A2(prog_data[13]), .B1(\mem[33][13] ), .B2(n7089), .Z(n4138) );
  OA22D0 U3599 ( .A1(n7090), .A2(prog_data[12]), .B1(\mem[33][12] ), .B2(n7089), .Z(n4137) );
  OA22D0 U3600 ( .A1(n7090), .A2(prog_data[11]), .B1(\mem[33][11] ), .B2(n7089), .Z(n4136) );
  OA22D0 U3601 ( .A1(n7090), .A2(prog_data[10]), .B1(\mem[33][10] ), .B2(n7089), .Z(n4135) );
  OA22D0 U3602 ( .A1(n7090), .A2(prog_data[9]), .B1(\mem[33][9] ), .B2(n7089), 
        .Z(n4134) );
  OA22D0 U3603 ( .A1(n7090), .A2(prog_data[8]), .B1(\mem[33][8] ), .B2(n7089), 
        .Z(n4133) );
  OA22D0 U3604 ( .A1(n7090), .A2(prog_data[7]), .B1(\mem[33][7] ), .B2(n7089), 
        .Z(n4132) );
  OA22D0 U3605 ( .A1(n7090), .A2(prog_data[6]), .B1(\mem[33][6] ), .B2(n7089), 
        .Z(n4131) );
  OA22D0 U3606 ( .A1(n7090), .A2(prog_data[5]), .B1(\mem[33][5] ), .B2(n7089), 
        .Z(n4130) );
  OA22D0 U3607 ( .A1(n7090), .A2(prog_data[4]), .B1(\mem[33][4] ), .B2(n7089), 
        .Z(n4129) );
  OA22D0 U3608 ( .A1(n7090), .A2(prog_data[3]), .B1(\mem[33][3] ), .B2(n7089), 
        .Z(n4128) );
  OA22D0 U3609 ( .A1(n7090), .A2(prog_data[2]), .B1(\mem[33][2] ), .B2(n7089), 
        .Z(n4127) );
  OA22D0 U3610 ( .A1(n7090), .A2(prog_data[1]), .B1(\mem[33][1] ), .B2(n7089), 
        .Z(n4126) );
  OA22D0 U3611 ( .A1(n7090), .A2(prog_data[0]), .B1(\mem[33][0] ), .B2(n7089), 
        .Z(n4125) );
  NR2D0 U3612 ( .A1(n7534), .A2(n7117), .ZN(n7091) );
  INVD0 U3613 ( .I(n7091), .ZN(n7092) );
  OA22D0 U3614 ( .A1(n7092), .A2(prog_data[15]), .B1(\mem[34][15] ), .B2(n7091), .Z(n4124) );
  OA22D0 U3615 ( .A1(n7092), .A2(prog_data[14]), .B1(\mem[34][14] ), .B2(n7091), .Z(n4123) );
  OA22D0 U3616 ( .A1(n7092), .A2(prog_data[13]), .B1(\mem[34][13] ), .B2(n7091), .Z(n4122) );
  OA22D0 U3617 ( .A1(n7092), .A2(prog_data[12]), .B1(\mem[34][12] ), .B2(n7091), .Z(n4121) );
  OA22D0 U3618 ( .A1(n7092), .A2(prog_data[11]), .B1(\mem[34][11] ), .B2(n7091), .Z(n4120) );
  OA22D0 U3619 ( .A1(n7092), .A2(prog_data[10]), .B1(\mem[34][10] ), .B2(n7091), .Z(n4119) );
  OA22D0 U3620 ( .A1(n7092), .A2(prog_data[9]), .B1(\mem[34][9] ), .B2(n7091), 
        .Z(n4118) );
  OA22D0 U3621 ( .A1(n7092), .A2(prog_data[8]), .B1(\mem[34][8] ), .B2(n7091), 
        .Z(n4117) );
  OA22D0 U3622 ( .A1(n7092), .A2(prog_data[7]), .B1(\mem[34][7] ), .B2(n7091), 
        .Z(n4116) );
  OA22D0 U3623 ( .A1(n7092), .A2(prog_data[6]), .B1(\mem[34][6] ), .B2(n7091), 
        .Z(n4115) );
  OA22D0 U3624 ( .A1(n7092), .A2(prog_data[5]), .B1(\mem[34][5] ), .B2(n7091), 
        .Z(n4114) );
  OA22D0 U3625 ( .A1(n7092), .A2(prog_data[4]), .B1(\mem[34][4] ), .B2(n7091), 
        .Z(n4113) );
  OA22D0 U3626 ( .A1(n7092), .A2(prog_data[3]), .B1(\mem[34][3] ), .B2(n7091), 
        .Z(n4112) );
  OA22D0 U3627 ( .A1(n7092), .A2(prog_data[2]), .B1(\mem[34][2] ), .B2(n7091), 
        .Z(n4111) );
  OA22D0 U3628 ( .A1(n7092), .A2(prog_data[1]), .B1(\mem[34][1] ), .B2(n7091), 
        .Z(n4110) );
  OA22D0 U3629 ( .A1(n7092), .A2(prog_data[0]), .B1(\mem[34][0] ), .B2(n7091), 
        .Z(n4109) );
  NR2D0 U3630 ( .A1(n7537), .A2(n7117), .ZN(n7093) );
  INVD0 U3631 ( .I(n7093), .ZN(n7094) );
  OA22D0 U3632 ( .A1(n7094), .A2(prog_data[15]), .B1(\mem[35][15] ), .B2(n7093), .Z(n4108) );
  OA22D0 U3633 ( .A1(n7094), .A2(prog_data[14]), .B1(\mem[35][14] ), .B2(n7093), .Z(n4107) );
  OA22D0 U3634 ( .A1(n7094), .A2(prog_data[13]), .B1(\mem[35][13] ), .B2(n7093), .Z(n4106) );
  OA22D0 U3635 ( .A1(n7094), .A2(prog_data[12]), .B1(\mem[35][12] ), .B2(n7093), .Z(n4105) );
  OA22D0 U3636 ( .A1(n7094), .A2(prog_data[11]), .B1(\mem[35][11] ), .B2(n7093), .Z(n4104) );
  OA22D0 U3637 ( .A1(n7094), .A2(prog_data[10]), .B1(\mem[35][10] ), .B2(n7093), .Z(n4103) );
  OA22D0 U3638 ( .A1(n7094), .A2(prog_data[9]), .B1(\mem[35][9] ), .B2(n7093), 
        .Z(n4102) );
  OA22D0 U3639 ( .A1(n7094), .A2(prog_data[8]), .B1(\mem[35][8] ), .B2(n7093), 
        .Z(n4101) );
  OA22D0 U3640 ( .A1(n7094), .A2(prog_data[7]), .B1(\mem[35][7] ), .B2(n7093), 
        .Z(n4100) );
  OA22D0 U3641 ( .A1(n7094), .A2(prog_data[6]), .B1(\mem[35][6] ), .B2(n7093), 
        .Z(n4099) );
  OA22D0 U3642 ( .A1(n7094), .A2(prog_data[5]), .B1(\mem[35][5] ), .B2(n7093), 
        .Z(n4098) );
  OA22D0 U3643 ( .A1(n7094), .A2(prog_data[4]), .B1(\mem[35][4] ), .B2(n7093), 
        .Z(n4097) );
  OA22D0 U3644 ( .A1(n7094), .A2(prog_data[3]), .B1(\mem[35][3] ), .B2(n7093), 
        .Z(n4096) );
  OA22D0 U3645 ( .A1(n7094), .A2(prog_data[2]), .B1(\mem[35][2] ), .B2(n7093), 
        .Z(n4095) );
  OA22D0 U3646 ( .A1(n7094), .A2(prog_data[1]), .B1(\mem[35][1] ), .B2(n7093), 
        .Z(n4094) );
  OA22D0 U3647 ( .A1(n7094), .A2(prog_data[0]), .B1(\mem[35][0] ), .B2(n7093), 
        .Z(n4093) );
  NR2D0 U3648 ( .A1(n7540), .A2(n7117), .ZN(n7095) );
  INVD0 U3649 ( .I(n7095), .ZN(n7096) );
  OA22D0 U3650 ( .A1(n7096), .A2(prog_data[15]), .B1(\mem[36][15] ), .B2(n7095), .Z(n4092) );
  OA22D0 U3651 ( .A1(n7096), .A2(prog_data[14]), .B1(\mem[36][14] ), .B2(n7095), .Z(n4091) );
  OA22D0 U3652 ( .A1(n7096), .A2(prog_data[13]), .B1(\mem[36][13] ), .B2(n7095), .Z(n4090) );
  OA22D0 U3653 ( .A1(n7096), .A2(prog_data[12]), .B1(\mem[36][12] ), .B2(n7095), .Z(n4089) );
  OA22D0 U3654 ( .A1(n7096), .A2(prog_data[11]), .B1(\mem[36][11] ), .B2(n7095), .Z(n4088) );
  OA22D0 U3655 ( .A1(n7096), .A2(prog_data[10]), .B1(\mem[36][10] ), .B2(n7095), .Z(n4087) );
  OA22D0 U3656 ( .A1(n7096), .A2(prog_data[9]), .B1(\mem[36][9] ), .B2(n7095), 
        .Z(n4086) );
  OA22D0 U3657 ( .A1(n7096), .A2(prog_data[8]), .B1(\mem[36][8] ), .B2(n7095), 
        .Z(n4085) );
  OA22D0 U3658 ( .A1(n7096), .A2(prog_data[7]), .B1(\mem[36][7] ), .B2(n7095), 
        .Z(n4084) );
  OA22D0 U3659 ( .A1(n7096), .A2(prog_data[6]), .B1(\mem[36][6] ), .B2(n7095), 
        .Z(n4083) );
  OA22D0 U3660 ( .A1(n7096), .A2(prog_data[5]), .B1(\mem[36][5] ), .B2(n7095), 
        .Z(n4082) );
  OA22D0 U3661 ( .A1(n7096), .A2(prog_data[4]), .B1(\mem[36][4] ), .B2(n7095), 
        .Z(n4081) );
  OA22D0 U3662 ( .A1(n7096), .A2(prog_data[3]), .B1(\mem[36][3] ), .B2(n7095), 
        .Z(n4080) );
  OA22D0 U3663 ( .A1(n7096), .A2(prog_data[2]), .B1(\mem[36][2] ), .B2(n7095), 
        .Z(n4079) );
  OA22D0 U3664 ( .A1(n7096), .A2(prog_data[1]), .B1(\mem[36][1] ), .B2(n7095), 
        .Z(n4078) );
  OA22D0 U3665 ( .A1(n7096), .A2(prog_data[0]), .B1(\mem[36][0] ), .B2(n7095), 
        .Z(n4077) );
  NR2D0 U3666 ( .A1(n7543), .A2(n7117), .ZN(n7097) );
  INVD0 U3667 ( .I(n7097), .ZN(n7098) );
  OA22D0 U3668 ( .A1(n7098), .A2(prog_data[15]), .B1(\mem[37][15] ), .B2(n7097), .Z(n4076) );
  OA22D0 U3669 ( .A1(n7098), .A2(prog_data[14]), .B1(\mem[37][14] ), .B2(n7097), .Z(n4075) );
  OA22D0 U3670 ( .A1(n7098), .A2(prog_data[13]), .B1(\mem[37][13] ), .B2(n7097), .Z(n4074) );
  OA22D0 U3671 ( .A1(n7098), .A2(prog_data[12]), .B1(\mem[37][12] ), .B2(n7097), .Z(n4073) );
  OA22D0 U3672 ( .A1(n7098), .A2(prog_data[11]), .B1(\mem[37][11] ), .B2(n7097), .Z(n4072) );
  OA22D0 U3673 ( .A1(n7098), .A2(prog_data[10]), .B1(\mem[37][10] ), .B2(n7097), .Z(n4071) );
  OA22D0 U3674 ( .A1(n7098), .A2(prog_data[9]), .B1(\mem[37][9] ), .B2(n7097), 
        .Z(n4070) );
  OA22D0 U3675 ( .A1(n7098), .A2(prog_data[8]), .B1(\mem[37][8] ), .B2(n7097), 
        .Z(n4069) );
  OA22D0 U3676 ( .A1(n7098), .A2(prog_data[7]), .B1(\mem[37][7] ), .B2(n7097), 
        .Z(n4068) );
  OA22D0 U3677 ( .A1(n7098), .A2(prog_data[6]), .B1(\mem[37][6] ), .B2(n7097), 
        .Z(n4067) );
  OA22D0 U3678 ( .A1(n7098), .A2(prog_data[5]), .B1(\mem[37][5] ), .B2(n7097), 
        .Z(n4066) );
  OA22D0 U3679 ( .A1(n7098), .A2(prog_data[4]), .B1(\mem[37][4] ), .B2(n7097), 
        .Z(n4065) );
  OA22D0 U3680 ( .A1(n7098), .A2(prog_data[3]), .B1(\mem[37][3] ), .B2(n7097), 
        .Z(n4064) );
  OA22D0 U3681 ( .A1(n7098), .A2(prog_data[2]), .B1(\mem[37][2] ), .B2(n7097), 
        .Z(n4063) );
  OA22D0 U3682 ( .A1(n7098), .A2(prog_data[1]), .B1(\mem[37][1] ), .B2(n7097), 
        .Z(n4062) );
  OA22D0 U3683 ( .A1(n7098), .A2(prog_data[0]), .B1(\mem[37][0] ), .B2(n7097), 
        .Z(n4061) );
  NR2D0 U3684 ( .A1(n7546), .A2(n7117), .ZN(n7099) );
  INVD0 U3685 ( .I(n7099), .ZN(n7100) );
  OA22D0 U3686 ( .A1(n7100), .A2(prog_data[15]), .B1(\mem[38][15] ), .B2(n7099), .Z(n4060) );
  OA22D0 U3687 ( .A1(n7100), .A2(prog_data[14]), .B1(\mem[38][14] ), .B2(n7099), .Z(n4059) );
  OA22D0 U3688 ( .A1(n7100), .A2(prog_data[13]), .B1(\mem[38][13] ), .B2(n7099), .Z(n4058) );
  OA22D0 U3689 ( .A1(n7100), .A2(prog_data[12]), .B1(\mem[38][12] ), .B2(n7099), .Z(n4057) );
  OA22D0 U3690 ( .A1(n7100), .A2(prog_data[11]), .B1(\mem[38][11] ), .B2(n7099), .Z(n4056) );
  OA22D0 U3691 ( .A1(n7100), .A2(prog_data[10]), .B1(\mem[38][10] ), .B2(n7099), .Z(n4055) );
  OA22D0 U3692 ( .A1(n7100), .A2(prog_data[9]), .B1(\mem[38][9] ), .B2(n7099), 
        .Z(n4054) );
  OA22D0 U3693 ( .A1(n7100), .A2(prog_data[8]), .B1(\mem[38][8] ), .B2(n7099), 
        .Z(n4053) );
  OA22D0 U3694 ( .A1(n7100), .A2(prog_data[7]), .B1(\mem[38][7] ), .B2(n7099), 
        .Z(n4052) );
  OA22D0 U3695 ( .A1(n7100), .A2(prog_data[6]), .B1(\mem[38][6] ), .B2(n7099), 
        .Z(n4051) );
  OA22D0 U3696 ( .A1(n7100), .A2(prog_data[5]), .B1(\mem[38][5] ), .B2(n7099), 
        .Z(n4050) );
  OA22D0 U3697 ( .A1(n7100), .A2(prog_data[4]), .B1(\mem[38][4] ), .B2(n7099), 
        .Z(n4049) );
  OA22D0 U3698 ( .A1(n7100), .A2(prog_data[3]), .B1(\mem[38][3] ), .B2(n7099), 
        .Z(n4048) );
  OA22D0 U3699 ( .A1(n7100), .A2(prog_data[2]), .B1(\mem[38][2] ), .B2(n7099), 
        .Z(n4047) );
  OA22D0 U3700 ( .A1(n7100), .A2(prog_data[1]), .B1(\mem[38][1] ), .B2(n7099), 
        .Z(n4046) );
  OA22D0 U3701 ( .A1(n7100), .A2(prog_data[0]), .B1(\mem[38][0] ), .B2(n7099), 
        .Z(n4045) );
  NR2D0 U3702 ( .A1(n7549), .A2(n7117), .ZN(n7101) );
  OA22D0 U3703 ( .A1(n7102), .A2(prog_data[15]), .B1(\mem[39][15] ), .B2(n7101), .Z(n4044) );
  OA22D0 U3704 ( .A1(n7102), .A2(prog_data[14]), .B1(\mem[39][14] ), .B2(n7101), .Z(n4043) );
  OA22D0 U3705 ( .A1(n7102), .A2(prog_data[13]), .B1(\mem[39][13] ), .B2(n7101), .Z(n4042) );
  OA22D0 U3706 ( .A1(n7102), .A2(prog_data[12]), .B1(\mem[39][12] ), .B2(n7101), .Z(n4041) );
  OA22D0 U3707 ( .A1(n7102), .A2(prog_data[11]), .B1(\mem[39][11] ), .B2(n7101), .Z(n4040) );
  OA22D0 U3708 ( .A1(n7102), .A2(prog_data[10]), .B1(\mem[39][10] ), .B2(n7101), .Z(n4039) );
  OA22D0 U3709 ( .A1(n7102), .A2(prog_data[9]), .B1(\mem[39][9] ), .B2(n7101), 
        .Z(n4038) );
  OA22D0 U3710 ( .A1(n7102), .A2(prog_data[8]), .B1(\mem[39][8] ), .B2(n7101), 
        .Z(n4037) );
  OA22D0 U3711 ( .A1(n7102), .A2(prog_data[7]), .B1(\mem[39][7] ), .B2(n7101), 
        .Z(n4036) );
  OA22D0 U3712 ( .A1(n7102), .A2(prog_data[6]), .B1(\mem[39][6] ), .B2(n7101), 
        .Z(n4035) );
  OA22D0 U3713 ( .A1(n7102), .A2(prog_data[5]), .B1(\mem[39][5] ), .B2(n7101), 
        .Z(n4034) );
  OA22D0 U3714 ( .A1(n7102), .A2(prog_data[4]), .B1(\mem[39][4] ), .B2(n7101), 
        .Z(n4033) );
  OA22D0 U3715 ( .A1(n7102), .A2(prog_data[3]), .B1(\mem[39][3] ), .B2(n7101), 
        .Z(n4032) );
  OA22D0 U3716 ( .A1(n7102), .A2(prog_data[2]), .B1(\mem[39][2] ), .B2(n7101), 
        .Z(n4031) );
  OA22D0 U3717 ( .A1(n7102), .A2(prog_data[1]), .B1(\mem[39][1] ), .B2(n7101), 
        .Z(n4030) );
  OA22D0 U3718 ( .A1(n7102), .A2(prog_data[0]), .B1(\mem[39][0] ), .B2(n7101), 
        .Z(n4029) );
  NR2D0 U3719 ( .A1(n7552), .A2(n7117), .ZN(n7103) );
  INVD0 U3720 ( .I(n7103), .ZN(n7104) );
  OA22D0 U3721 ( .A1(n7104), .A2(prog_data[15]), .B1(\mem[40][15] ), .B2(n7103), .Z(n4028) );
  OA22D0 U3722 ( .A1(n7104), .A2(prog_data[14]), .B1(\mem[40][14] ), .B2(n7103), .Z(n4027) );
  OA22D0 U3723 ( .A1(n7104), .A2(prog_data[13]), .B1(\mem[40][13] ), .B2(n7103), .Z(n4026) );
  OA22D0 U3724 ( .A1(n7104), .A2(prog_data[12]), .B1(\mem[40][12] ), .B2(n7103), .Z(n4025) );
  OA22D0 U3725 ( .A1(n7104), .A2(prog_data[11]), .B1(\mem[40][11] ), .B2(n7103), .Z(n4024) );
  OA22D0 U3726 ( .A1(n7104), .A2(prog_data[10]), .B1(\mem[40][10] ), .B2(n7103), .Z(n4023) );
  OA22D0 U3727 ( .A1(n7104), .A2(prog_data[9]), .B1(\mem[40][9] ), .B2(n7103), 
        .Z(n4022) );
  OA22D0 U3728 ( .A1(n7104), .A2(prog_data[8]), .B1(\mem[40][8] ), .B2(n7103), 
        .Z(n4021) );
  OA22D0 U3729 ( .A1(n7104), .A2(prog_data[7]), .B1(\mem[40][7] ), .B2(n7103), 
        .Z(n4020) );
  OA22D0 U3730 ( .A1(n7104), .A2(prog_data[6]), .B1(\mem[40][6] ), .B2(n7103), 
        .Z(n4019) );
  OA22D0 U3731 ( .A1(n7104), .A2(prog_data[5]), .B1(\mem[40][5] ), .B2(n7103), 
        .Z(n4018) );
  OA22D0 U3732 ( .A1(n7104), .A2(prog_data[4]), .B1(\mem[40][4] ), .B2(n7103), 
        .Z(n4017) );
  OA22D0 U3733 ( .A1(n7104), .A2(prog_data[3]), .B1(\mem[40][3] ), .B2(n7103), 
        .Z(n4016) );
  OA22D0 U3734 ( .A1(n7104), .A2(prog_data[2]), .B1(\mem[40][2] ), .B2(n7103), 
        .Z(n4015) );
  OA22D0 U3735 ( .A1(n7104), .A2(prog_data[1]), .B1(\mem[40][1] ), .B2(n7103), 
        .Z(n4014) );
  OA22D0 U3736 ( .A1(n7104), .A2(prog_data[0]), .B1(\mem[40][0] ), .B2(n7103), 
        .Z(n4013) );
  NR2D0 U3737 ( .A1(n7555), .A2(n7117), .ZN(n7105) );
  INVD0 U3738 ( .I(n7105), .ZN(n7106) );
  OA22D0 U3739 ( .A1(n7106), .A2(prog_data[15]), .B1(\mem[41][15] ), .B2(n7105), .Z(n4012) );
  OA22D0 U3740 ( .A1(n7106), .A2(prog_data[14]), .B1(\mem[41][14] ), .B2(n7105), .Z(n4011) );
  OA22D0 U3741 ( .A1(n7106), .A2(prog_data[13]), .B1(\mem[41][13] ), .B2(n7105), .Z(n4010) );
  OA22D0 U3742 ( .A1(n7106), .A2(prog_data[12]), .B1(\mem[41][12] ), .B2(n7105), .Z(n4009) );
  OA22D0 U3743 ( .A1(n7106), .A2(prog_data[11]), .B1(\mem[41][11] ), .B2(n7105), .Z(n4008) );
  OA22D0 U3744 ( .A1(n7106), .A2(prog_data[10]), .B1(\mem[41][10] ), .B2(n7105), .Z(n4007) );
  OA22D0 U3745 ( .A1(n7106), .A2(prog_data[9]), .B1(\mem[41][9] ), .B2(n7105), 
        .Z(n4006) );
  OA22D0 U3746 ( .A1(n7106), .A2(prog_data[8]), .B1(\mem[41][8] ), .B2(n7105), 
        .Z(n4005) );
  OA22D0 U3747 ( .A1(n7106), .A2(prog_data[7]), .B1(\mem[41][7] ), .B2(n7105), 
        .Z(n4004) );
  OA22D0 U3748 ( .A1(n7106), .A2(prog_data[6]), .B1(\mem[41][6] ), .B2(n7105), 
        .Z(n4003) );
  OA22D0 U3749 ( .A1(n7106), .A2(prog_data[5]), .B1(\mem[41][5] ), .B2(n7105), 
        .Z(n4002) );
  OA22D0 U3750 ( .A1(n7106), .A2(prog_data[4]), .B1(\mem[41][4] ), .B2(n7105), 
        .Z(n4001) );
  OA22D0 U3751 ( .A1(n7106), .A2(prog_data[3]), .B1(\mem[41][3] ), .B2(n7105), 
        .Z(n4000) );
  OA22D0 U3752 ( .A1(n7106), .A2(prog_data[2]), .B1(\mem[41][2] ), .B2(n7105), 
        .Z(n3999) );
  OA22D0 U3753 ( .A1(n7106), .A2(prog_data[1]), .B1(\mem[41][1] ), .B2(n7105), 
        .Z(n3998) );
  OA22D0 U3754 ( .A1(n7106), .A2(prog_data[0]), .B1(\mem[41][0] ), .B2(n7105), 
        .Z(n3997) );
  NR2D0 U3755 ( .A1(n7558), .A2(n7117), .ZN(n7107) );
  INVD0 U3756 ( .I(n7107), .ZN(n7108) );
  OA22D0 U3757 ( .A1(n7108), .A2(prog_data[15]), .B1(\mem[42][15] ), .B2(n7107), .Z(n3996) );
  OA22D0 U3758 ( .A1(n7108), .A2(prog_data[14]), .B1(\mem[42][14] ), .B2(n7107), .Z(n3995) );
  OA22D0 U3759 ( .A1(n7108), .A2(prog_data[13]), .B1(\mem[42][13] ), .B2(n7107), .Z(n3994) );
  OA22D0 U3760 ( .A1(n7108), .A2(prog_data[12]), .B1(\mem[42][12] ), .B2(n7107), .Z(n3993) );
  OA22D0 U3761 ( .A1(n7108), .A2(prog_data[11]), .B1(\mem[42][11] ), .B2(n7107), .Z(n3992) );
  OA22D0 U3762 ( .A1(n7108), .A2(prog_data[10]), .B1(\mem[42][10] ), .B2(n7107), .Z(n3991) );
  OA22D0 U3763 ( .A1(n7108), .A2(prog_data[9]), .B1(\mem[42][9] ), .B2(n7107), 
        .Z(n3990) );
  OA22D0 U3764 ( .A1(n7108), .A2(prog_data[8]), .B1(\mem[42][8] ), .B2(n7107), 
        .Z(n3989) );
  OA22D0 U3765 ( .A1(n7108), .A2(prog_data[7]), .B1(\mem[42][7] ), .B2(n7107), 
        .Z(n3988) );
  OA22D0 U3766 ( .A1(n7108), .A2(prog_data[6]), .B1(\mem[42][6] ), .B2(n7107), 
        .Z(n3987) );
  OA22D0 U3767 ( .A1(n7108), .A2(prog_data[5]), .B1(\mem[42][5] ), .B2(n7107), 
        .Z(n3986) );
  OA22D0 U3768 ( .A1(n7108), .A2(prog_data[4]), .B1(\mem[42][4] ), .B2(n7107), 
        .Z(n3985) );
  OA22D0 U3769 ( .A1(n7108), .A2(prog_data[3]), .B1(\mem[42][3] ), .B2(n7107), 
        .Z(n3984) );
  OA22D0 U3770 ( .A1(n7108), .A2(prog_data[2]), .B1(\mem[42][2] ), .B2(n7107), 
        .Z(n3983) );
  OA22D0 U3771 ( .A1(n7108), .A2(prog_data[1]), .B1(\mem[42][1] ), .B2(n7107), 
        .Z(n3982) );
  OA22D0 U3772 ( .A1(n7108), .A2(prog_data[0]), .B1(\mem[42][0] ), .B2(n7107), 
        .Z(n3981) );
  NR2D0 U3773 ( .A1(n7561), .A2(n7117), .ZN(n7109) );
  INVD0 U3774 ( .I(n7109), .ZN(n7110) );
  OA22D0 U3775 ( .A1(n7110), .A2(prog_data[15]), .B1(\mem[43][15] ), .B2(n7109), .Z(n3980) );
  OA22D0 U3776 ( .A1(n7110), .A2(prog_data[14]), .B1(\mem[43][14] ), .B2(n7109), .Z(n3979) );
  OA22D0 U3777 ( .A1(n7110), .A2(prog_data[13]), .B1(\mem[43][13] ), .B2(n7109), .Z(n3978) );
  OA22D0 U3778 ( .A1(n7110), .A2(prog_data[12]), .B1(\mem[43][12] ), .B2(n7109), .Z(n3977) );
  OA22D0 U3779 ( .A1(n7110), .A2(prog_data[11]), .B1(\mem[43][11] ), .B2(n7109), .Z(n3976) );
  OA22D0 U3780 ( .A1(n7110), .A2(prog_data[10]), .B1(\mem[43][10] ), .B2(n7109), .Z(n3975) );
  OA22D0 U3781 ( .A1(n7110), .A2(prog_data[9]), .B1(\mem[43][9] ), .B2(n7109), 
        .Z(n3974) );
  OA22D0 U3782 ( .A1(n7110), .A2(prog_data[8]), .B1(\mem[43][8] ), .B2(n7109), 
        .Z(n3973) );
  OA22D0 U3783 ( .A1(n7110), .A2(prog_data[7]), .B1(\mem[43][7] ), .B2(n7109), 
        .Z(n3972) );
  OA22D0 U3784 ( .A1(n7110), .A2(prog_data[6]), .B1(\mem[43][6] ), .B2(n7109), 
        .Z(n3971) );
  OA22D0 U3785 ( .A1(n7110), .A2(prog_data[5]), .B1(\mem[43][5] ), .B2(n7109), 
        .Z(n3970) );
  OA22D0 U3786 ( .A1(n7110), .A2(prog_data[4]), .B1(\mem[43][4] ), .B2(n7109), 
        .Z(n3969) );
  OA22D0 U3787 ( .A1(n7110), .A2(prog_data[3]), .B1(\mem[43][3] ), .B2(n7109), 
        .Z(n3968) );
  OA22D0 U3788 ( .A1(n7110), .A2(prog_data[2]), .B1(\mem[43][2] ), .B2(n7109), 
        .Z(n3967) );
  OA22D0 U3789 ( .A1(n7110), .A2(prog_data[1]), .B1(\mem[43][1] ), .B2(n7109), 
        .Z(n3966) );
  OA22D0 U3790 ( .A1(n7110), .A2(prog_data[0]), .B1(\mem[43][0] ), .B2(n7109), 
        .Z(n3965) );
  NR2D0 U3791 ( .A1(n7564), .A2(n7117), .ZN(n7111) );
  INVD0 U3792 ( .I(n7111), .ZN(n7112) );
  OA22D0 U3793 ( .A1(n7112), .A2(prog_data[15]), .B1(\mem[44][15] ), .B2(n7111), .Z(n3964) );
  OA22D0 U3794 ( .A1(n7112), .A2(prog_data[14]), .B1(\mem[44][14] ), .B2(n7111), .Z(n3963) );
  OA22D0 U3795 ( .A1(n7112), .A2(prog_data[13]), .B1(\mem[44][13] ), .B2(n7111), .Z(n3962) );
  OA22D0 U3796 ( .A1(n7112), .A2(prog_data[12]), .B1(\mem[44][12] ), .B2(n7111), .Z(n3961) );
  OA22D0 U3797 ( .A1(n7112), .A2(prog_data[11]), .B1(\mem[44][11] ), .B2(n7111), .Z(n3960) );
  OA22D0 U3798 ( .A1(n7112), .A2(prog_data[10]), .B1(\mem[44][10] ), .B2(n7111), .Z(n3959) );
  OA22D0 U3799 ( .A1(n7112), .A2(prog_data[9]), .B1(\mem[44][9] ), .B2(n7111), 
        .Z(n3958) );
  OA22D0 U3800 ( .A1(n7112), .A2(prog_data[8]), .B1(\mem[44][8] ), .B2(n7111), 
        .Z(n3957) );
  OA22D0 U3801 ( .A1(n7112), .A2(prog_data[7]), .B1(\mem[44][7] ), .B2(n7111), 
        .Z(n3956) );
  OA22D0 U3802 ( .A1(n7112), .A2(prog_data[6]), .B1(\mem[44][6] ), .B2(n7111), 
        .Z(n3955) );
  OA22D0 U3803 ( .A1(n7112), .A2(prog_data[5]), .B1(\mem[44][5] ), .B2(n7111), 
        .Z(n3954) );
  OA22D0 U3804 ( .A1(n7112), .A2(prog_data[4]), .B1(\mem[44][4] ), .B2(n7111), 
        .Z(n3953) );
  OA22D0 U3805 ( .A1(n7112), .A2(prog_data[3]), .B1(\mem[44][3] ), .B2(n7111), 
        .Z(n3952) );
  OA22D0 U3806 ( .A1(n7112), .A2(prog_data[2]), .B1(\mem[44][2] ), .B2(n7111), 
        .Z(n3951) );
  OA22D0 U3807 ( .A1(n7112), .A2(prog_data[1]), .B1(\mem[44][1] ), .B2(n7111), 
        .Z(n3950) );
  OA22D0 U3808 ( .A1(n7112), .A2(prog_data[0]), .B1(\mem[44][0] ), .B2(n7111), 
        .Z(n3949) );
  NR2D0 U3809 ( .A1(n7567), .A2(n7117), .ZN(n7113) );
  INVD0 U3810 ( .I(n7113), .ZN(n7114) );
  OA22D0 U3811 ( .A1(n7114), .A2(prog_data[15]), .B1(\mem[45][15] ), .B2(n7113), .Z(n3948) );
  OA22D0 U3812 ( .A1(n7114), .A2(prog_data[14]), .B1(\mem[45][14] ), .B2(n7113), .Z(n3947) );
  OA22D0 U3813 ( .A1(n7114), .A2(prog_data[13]), .B1(\mem[45][13] ), .B2(n7113), .Z(n3946) );
  OA22D0 U3814 ( .A1(n7114), .A2(prog_data[12]), .B1(\mem[45][12] ), .B2(n7113), .Z(n3945) );
  OA22D0 U3815 ( .A1(n7114), .A2(prog_data[11]), .B1(\mem[45][11] ), .B2(n7113), .Z(n3944) );
  OA22D0 U3816 ( .A1(n7114), .A2(prog_data[10]), .B1(\mem[45][10] ), .B2(n7113), .Z(n3943) );
  OA22D0 U3817 ( .A1(n7114), .A2(prog_data[9]), .B1(\mem[45][9] ), .B2(n7113), 
        .Z(n3942) );
  OA22D0 U3818 ( .A1(n7114), .A2(prog_data[8]), .B1(\mem[45][8] ), .B2(n7113), 
        .Z(n3941) );
  OA22D0 U3819 ( .A1(n7114), .A2(prog_data[7]), .B1(\mem[45][7] ), .B2(n7113), 
        .Z(n3940) );
  OA22D0 U3820 ( .A1(n7114), .A2(prog_data[6]), .B1(\mem[45][6] ), .B2(n7113), 
        .Z(n3939) );
  OA22D0 U3821 ( .A1(n7114), .A2(prog_data[5]), .B1(\mem[45][5] ), .B2(n7113), 
        .Z(n3938) );
  OA22D0 U3822 ( .A1(n7114), .A2(prog_data[4]), .B1(\mem[45][4] ), .B2(n7113), 
        .Z(n3937) );
  OA22D0 U3823 ( .A1(n7114), .A2(prog_data[3]), .B1(\mem[45][3] ), .B2(n7113), 
        .Z(n3936) );
  OA22D0 U3824 ( .A1(n7114), .A2(prog_data[2]), .B1(\mem[45][2] ), .B2(n7113), 
        .Z(n3935) );
  OA22D0 U3825 ( .A1(n7114), .A2(prog_data[1]), .B1(\mem[45][1] ), .B2(n7113), 
        .Z(n3934) );
  OA22D0 U3826 ( .A1(n7114), .A2(prog_data[0]), .B1(\mem[45][0] ), .B2(n7113), 
        .Z(n3933) );
  INVD0 U3827 ( .I(n7115), .ZN(n7116) );
  OA22D0 U3828 ( .A1(n7116), .A2(prog_data[15]), .B1(\mem[46][15] ), .B2(n7115), .Z(n3932) );
  OA22D0 U3829 ( .A1(n7116), .A2(prog_data[14]), .B1(\mem[46][14] ), .B2(n7115), .Z(n3931) );
  OA22D0 U3830 ( .A1(n7116), .A2(prog_data[13]), .B1(\mem[46][13] ), .B2(n7115), .Z(n3930) );
  OA22D0 U3831 ( .A1(n7116), .A2(prog_data[12]), .B1(\mem[46][12] ), .B2(n7115), .Z(n3929) );
  OA22D0 U3832 ( .A1(n7116), .A2(prog_data[11]), .B1(\mem[46][11] ), .B2(n7115), .Z(n3928) );
  OA22D0 U3833 ( .A1(n7116), .A2(prog_data[10]), .B1(\mem[46][10] ), .B2(n7115), .Z(n3927) );
  OA22D0 U3834 ( .A1(n7116), .A2(prog_data[9]), .B1(\mem[46][9] ), .B2(n7115), 
        .Z(n3926) );
  OA22D0 U3835 ( .A1(n7116), .A2(prog_data[8]), .B1(\mem[46][8] ), .B2(n7115), 
        .Z(n3925) );
  OA22D0 U3836 ( .A1(n7116), .A2(prog_data[7]), .B1(\mem[46][7] ), .B2(n7115), 
        .Z(n3924) );
  OA22D0 U3837 ( .A1(n7116), .A2(prog_data[6]), .B1(\mem[46][6] ), .B2(n7115), 
        .Z(n3923) );
  OA22D0 U3838 ( .A1(n7116), .A2(prog_data[5]), .B1(\mem[46][5] ), .B2(n7115), 
        .Z(n3922) );
  OA22D0 U3839 ( .A1(n7116), .A2(prog_data[4]), .B1(\mem[46][4] ), .B2(n7115), 
        .Z(n3921) );
  OA22D0 U3840 ( .A1(n7116), .A2(prog_data[3]), .B1(\mem[46][3] ), .B2(n7115), 
        .Z(n3920) );
  OA22D0 U3841 ( .A1(n7116), .A2(prog_data[2]), .B1(\mem[46][2] ), .B2(n7115), 
        .Z(n3919) );
  OA22D0 U3842 ( .A1(n7116), .A2(prog_data[1]), .B1(\mem[46][1] ), .B2(n7115), 
        .Z(n3918) );
  OA22D0 U3843 ( .A1(n7116), .A2(prog_data[0]), .B1(\mem[46][0] ), .B2(n7115), 
        .Z(n3917) );
  NR2D0 U3844 ( .A1(n7574), .A2(n7117), .ZN(n7118) );
  INVD0 U3845 ( .I(n7118), .ZN(n7119) );
  OA22D0 U3846 ( .A1(n7119), .A2(prog_data[15]), .B1(\mem[47][15] ), .B2(n7118), .Z(n3916) );
  OA22D0 U3847 ( .A1(n7119), .A2(prog_data[14]), .B1(\mem[47][14] ), .B2(n7118), .Z(n3915) );
  OA22D0 U3848 ( .A1(n7119), .A2(prog_data[13]), .B1(\mem[47][13] ), .B2(n7118), .Z(n3914) );
  OA22D0 U3849 ( .A1(n7119), .A2(prog_data[12]), .B1(\mem[47][12] ), .B2(n7118), .Z(n3913) );
  OA22D0 U3850 ( .A1(n7119), .A2(prog_data[11]), .B1(\mem[47][11] ), .B2(n7118), .Z(n3912) );
  OA22D0 U3851 ( .A1(n7119), .A2(prog_data[10]), .B1(\mem[47][10] ), .B2(n7118), .Z(n3911) );
  OA22D0 U3852 ( .A1(n7119), .A2(prog_data[9]), .B1(\mem[47][9] ), .B2(n7118), 
        .Z(n3910) );
  OA22D0 U3853 ( .A1(n7119), .A2(prog_data[8]), .B1(\mem[47][8] ), .B2(n7118), 
        .Z(n3909) );
  OA22D0 U3854 ( .A1(n7119), .A2(prog_data[7]), .B1(\mem[47][7] ), .B2(n7118), 
        .Z(n3908) );
  OA22D0 U3855 ( .A1(n7119), .A2(prog_data[6]), .B1(\mem[47][6] ), .B2(n7118), 
        .Z(n3907) );
  OA22D0 U3856 ( .A1(n7119), .A2(prog_data[5]), .B1(\mem[47][5] ), .B2(n7118), 
        .Z(n3906) );
  OA22D0 U3857 ( .A1(n7119), .A2(prog_data[4]), .B1(\mem[47][4] ), .B2(n7118), 
        .Z(n3905) );
  OA22D0 U3858 ( .A1(n7119), .A2(prog_data[3]), .B1(\mem[47][3] ), .B2(n7118), 
        .Z(n3904) );
  OA22D0 U3859 ( .A1(n7119), .A2(prog_data[2]), .B1(\mem[47][2] ), .B2(n7118), 
        .Z(n3903) );
  OA22D0 U3860 ( .A1(n7119), .A2(prog_data[1]), .B1(\mem[47][1] ), .B2(n7118), 
        .Z(n3902) );
  OA22D0 U3861 ( .A1(n7119), .A2(prog_data[0]), .B1(\mem[47][0] ), .B2(n7118), 
        .Z(n3901) );
  NR2D0 U3862 ( .A1(n7528), .A2(n7151), .ZN(n7121) );
  INVD0 U3863 ( .I(n7121), .ZN(n7122) );
  OA22D0 U3864 ( .A1(n7122), .A2(prog_data[15]), .B1(\mem[48][15] ), .B2(n7121), .Z(n3900) );
  OA22D0 U3865 ( .A1(n7122), .A2(prog_data[14]), .B1(\mem[48][14] ), .B2(n7121), .Z(n3899) );
  OA22D0 U3866 ( .A1(n7122), .A2(prog_data[13]), .B1(\mem[48][13] ), .B2(n7121), .Z(n3898) );
  OA22D0 U3867 ( .A1(n7122), .A2(prog_data[12]), .B1(\mem[48][12] ), .B2(n7121), .Z(n3897) );
  OA22D0 U3868 ( .A1(n7122), .A2(prog_data[11]), .B1(\mem[48][11] ), .B2(n7121), .Z(n3896) );
  OA22D0 U3869 ( .A1(n7122), .A2(prog_data[10]), .B1(\mem[48][10] ), .B2(n7121), .Z(n3895) );
  OA22D0 U3870 ( .A1(n7122), .A2(prog_data[9]), .B1(\mem[48][9] ), .B2(n7121), 
        .Z(n3894) );
  OA22D0 U3871 ( .A1(n7122), .A2(prog_data[8]), .B1(\mem[48][8] ), .B2(n7121), 
        .Z(n3893) );
  OA22D0 U3872 ( .A1(n7122), .A2(prog_data[7]), .B1(\mem[48][7] ), .B2(n7121), 
        .Z(n3892) );
  OA22D0 U3873 ( .A1(n7122), .A2(prog_data[6]), .B1(\mem[48][6] ), .B2(n7121), 
        .Z(n3891) );
  OA22D0 U3874 ( .A1(n7122), .A2(prog_data[5]), .B1(\mem[48][5] ), .B2(n7121), 
        .Z(n3890) );
  OA22D0 U3875 ( .A1(n7122), .A2(prog_data[4]), .B1(\mem[48][4] ), .B2(n7121), 
        .Z(n3889) );
  OA22D0 U3876 ( .A1(n7122), .A2(prog_data[3]), .B1(\mem[48][3] ), .B2(n7121), 
        .Z(n3888) );
  OA22D0 U3877 ( .A1(n7122), .A2(prog_data[2]), .B1(\mem[48][2] ), .B2(n7121), 
        .Z(n3887) );
  OA22D0 U3878 ( .A1(n7122), .A2(prog_data[1]), .B1(\mem[48][1] ), .B2(n7121), 
        .Z(n3886) );
  OA22D0 U3879 ( .A1(n7122), .A2(prog_data[0]), .B1(\mem[48][0] ), .B2(n7121), 
        .Z(n3885) );
  NR2D0 U3880 ( .A1(n7531), .A2(n7151), .ZN(n7123) );
  INVD0 U3881 ( .I(n7123), .ZN(n7124) );
  OA22D0 U3882 ( .A1(n7124), .A2(prog_data[15]), .B1(\mem[49][15] ), .B2(n7123), .Z(n3884) );
  OA22D0 U3883 ( .A1(n7124), .A2(prog_data[14]), .B1(\mem[49][14] ), .B2(n7123), .Z(n3883) );
  OA22D0 U3884 ( .A1(n7124), .A2(prog_data[13]), .B1(\mem[49][13] ), .B2(n7123), .Z(n3882) );
  OA22D0 U3885 ( .A1(n7124), .A2(prog_data[12]), .B1(\mem[49][12] ), .B2(n7123), .Z(n3881) );
  OA22D0 U3886 ( .A1(n7124), .A2(prog_data[11]), .B1(\mem[49][11] ), .B2(n7123), .Z(n3880) );
  OA22D0 U3887 ( .A1(n7124), .A2(prog_data[10]), .B1(\mem[49][10] ), .B2(n7123), .Z(n3879) );
  OA22D0 U3888 ( .A1(n7124), .A2(prog_data[9]), .B1(\mem[49][9] ), .B2(n7123), 
        .Z(n3878) );
  OA22D0 U3889 ( .A1(n7124), .A2(prog_data[8]), .B1(\mem[49][8] ), .B2(n7123), 
        .Z(n3877) );
  OA22D0 U3890 ( .A1(n7124), .A2(prog_data[7]), .B1(\mem[49][7] ), .B2(n7123), 
        .Z(n3876) );
  OA22D0 U3891 ( .A1(n7124), .A2(prog_data[6]), .B1(\mem[49][6] ), .B2(n7123), 
        .Z(n3875) );
  OA22D0 U3892 ( .A1(n7124), .A2(prog_data[5]), .B1(\mem[49][5] ), .B2(n7123), 
        .Z(n3874) );
  OA22D0 U3893 ( .A1(n7124), .A2(prog_data[4]), .B1(\mem[49][4] ), .B2(n7123), 
        .Z(n3873) );
  OA22D0 U3894 ( .A1(n7124), .A2(prog_data[3]), .B1(\mem[49][3] ), .B2(n7123), 
        .Z(n3872) );
  OA22D0 U3895 ( .A1(n7124), .A2(prog_data[2]), .B1(\mem[49][2] ), .B2(n7123), 
        .Z(n3871) );
  OA22D0 U3896 ( .A1(n7124), .A2(prog_data[1]), .B1(\mem[49][1] ), .B2(n7123), 
        .Z(n3870) );
  OA22D0 U3897 ( .A1(n7124), .A2(prog_data[0]), .B1(\mem[49][0] ), .B2(n7123), 
        .Z(n3869) );
  NR2D0 U3898 ( .A1(n7534), .A2(n7151), .ZN(n7125) );
  INVD0 U3899 ( .I(n7125), .ZN(n7126) );
  OA22D0 U3900 ( .A1(n7126), .A2(prog_data[15]), .B1(\mem[50][15] ), .B2(n7125), .Z(n3868) );
  OA22D0 U3901 ( .A1(n7126), .A2(prog_data[14]), .B1(\mem[50][14] ), .B2(n7125), .Z(n3867) );
  OA22D0 U3902 ( .A1(n7126), .A2(prog_data[13]), .B1(\mem[50][13] ), .B2(n7125), .Z(n3866) );
  OA22D0 U3903 ( .A1(n7126), .A2(prog_data[12]), .B1(\mem[50][12] ), .B2(n7125), .Z(n3865) );
  OA22D0 U3904 ( .A1(n7126), .A2(prog_data[11]), .B1(\mem[50][11] ), .B2(n7125), .Z(n3864) );
  OA22D0 U3905 ( .A1(n7126), .A2(prog_data[10]), .B1(\mem[50][10] ), .B2(n7125), .Z(n3863) );
  OA22D0 U3906 ( .A1(n7126), .A2(prog_data[9]), .B1(\mem[50][9] ), .B2(n7125), 
        .Z(n3862) );
  OA22D0 U3907 ( .A1(n7126), .A2(prog_data[8]), .B1(\mem[50][8] ), .B2(n7125), 
        .Z(n3861) );
  OA22D0 U3908 ( .A1(n7126), .A2(prog_data[7]), .B1(\mem[50][7] ), .B2(n7125), 
        .Z(n3860) );
  OA22D0 U3909 ( .A1(n7126), .A2(prog_data[6]), .B1(\mem[50][6] ), .B2(n7125), 
        .Z(n3859) );
  OA22D0 U3910 ( .A1(n7126), .A2(prog_data[5]), .B1(\mem[50][5] ), .B2(n7125), 
        .Z(n3858) );
  OA22D0 U3911 ( .A1(n7126), .A2(prog_data[4]), .B1(\mem[50][4] ), .B2(n7125), 
        .Z(n3857) );
  OA22D0 U3912 ( .A1(n7126), .A2(prog_data[3]), .B1(\mem[50][3] ), .B2(n7125), 
        .Z(n3856) );
  OA22D0 U3913 ( .A1(n7126), .A2(prog_data[2]), .B1(\mem[50][2] ), .B2(n7125), 
        .Z(n3855) );
  OA22D0 U3914 ( .A1(n7126), .A2(prog_data[1]), .B1(\mem[50][1] ), .B2(n7125), 
        .Z(n3854) );
  OA22D0 U3915 ( .A1(n7126), .A2(prog_data[0]), .B1(\mem[50][0] ), .B2(n7125), 
        .Z(n3853) );
  NR2D0 U3916 ( .A1(n7537), .A2(n7151), .ZN(n7127) );
  INVD0 U3917 ( .I(n7127), .ZN(n7128) );
  OA22D0 U3918 ( .A1(n7128), .A2(prog_data[15]), .B1(\mem[51][15] ), .B2(n7127), .Z(n3852) );
  OA22D0 U3919 ( .A1(n7128), .A2(prog_data[14]), .B1(\mem[51][14] ), .B2(n7127), .Z(n3851) );
  OA22D0 U3920 ( .A1(n7128), .A2(prog_data[13]), .B1(\mem[51][13] ), .B2(n7127), .Z(n3850) );
  OA22D0 U3921 ( .A1(n7128), .A2(prog_data[12]), .B1(\mem[51][12] ), .B2(n7127), .Z(n3849) );
  OA22D0 U3922 ( .A1(n7128), .A2(prog_data[11]), .B1(\mem[51][11] ), .B2(n7127), .Z(n3848) );
  OA22D0 U3923 ( .A1(n7128), .A2(prog_data[10]), .B1(\mem[51][10] ), .B2(n7127), .Z(n3847) );
  OA22D0 U3924 ( .A1(n7128), .A2(prog_data[9]), .B1(\mem[51][9] ), .B2(n7127), 
        .Z(n3846) );
  OA22D0 U3925 ( .A1(n7128), .A2(prog_data[8]), .B1(\mem[51][8] ), .B2(n7127), 
        .Z(n3845) );
  OA22D0 U3926 ( .A1(n7128), .A2(prog_data[7]), .B1(\mem[51][7] ), .B2(n7127), 
        .Z(n3844) );
  OA22D0 U3927 ( .A1(n7128), .A2(prog_data[6]), .B1(\mem[51][6] ), .B2(n7127), 
        .Z(n3843) );
  OA22D0 U3928 ( .A1(n7128), .A2(prog_data[5]), .B1(\mem[51][5] ), .B2(n7127), 
        .Z(n3842) );
  OA22D0 U3929 ( .A1(n7128), .A2(prog_data[4]), .B1(\mem[51][4] ), .B2(n7127), 
        .Z(n3841) );
  OA22D0 U3930 ( .A1(n7128), .A2(prog_data[3]), .B1(\mem[51][3] ), .B2(n7127), 
        .Z(n3840) );
  OA22D0 U3931 ( .A1(n7128), .A2(prog_data[2]), .B1(\mem[51][2] ), .B2(n7127), 
        .Z(n3839) );
  OA22D0 U3932 ( .A1(n7128), .A2(prog_data[1]), .B1(\mem[51][1] ), .B2(n7127), 
        .Z(n3838) );
  OA22D0 U3933 ( .A1(n7128), .A2(prog_data[0]), .B1(\mem[51][0] ), .B2(n7127), 
        .Z(n3837) );
  NR2D0 U3934 ( .A1(n7540), .A2(n7151), .ZN(n7129) );
  INVD0 U3935 ( .I(n7129), .ZN(n7130) );
  OA22D0 U3936 ( .A1(n7130), .A2(prog_data[15]), .B1(\mem[52][15] ), .B2(n7129), .Z(n3836) );
  OA22D0 U3937 ( .A1(n7130), .A2(prog_data[14]), .B1(\mem[52][14] ), .B2(n7129), .Z(n3835) );
  OA22D0 U3938 ( .A1(n7130), .A2(prog_data[13]), .B1(\mem[52][13] ), .B2(n7129), .Z(n3834) );
  OA22D0 U3939 ( .A1(n7130), .A2(prog_data[12]), .B1(\mem[52][12] ), .B2(n7129), .Z(n3833) );
  OA22D0 U3940 ( .A1(n7130), .A2(prog_data[11]), .B1(\mem[52][11] ), .B2(n7129), .Z(n3832) );
  OA22D0 U3941 ( .A1(n7130), .A2(prog_data[10]), .B1(\mem[52][10] ), .B2(n7129), .Z(n3831) );
  OA22D0 U3942 ( .A1(n7130), .A2(prog_data[9]), .B1(\mem[52][9] ), .B2(n7129), 
        .Z(n3830) );
  OA22D0 U3943 ( .A1(n7130), .A2(prog_data[8]), .B1(\mem[52][8] ), .B2(n7129), 
        .Z(n3829) );
  OA22D0 U3944 ( .A1(n7130), .A2(prog_data[7]), .B1(\mem[52][7] ), .B2(n7129), 
        .Z(n3828) );
  OA22D0 U3945 ( .A1(n7130), .A2(prog_data[6]), .B1(\mem[52][6] ), .B2(n7129), 
        .Z(n3827) );
  OA22D0 U3946 ( .A1(n7130), .A2(prog_data[5]), .B1(\mem[52][5] ), .B2(n7129), 
        .Z(n3826) );
  OA22D0 U3947 ( .A1(n7130), .A2(prog_data[4]), .B1(\mem[52][4] ), .B2(n7129), 
        .Z(n3825) );
  OA22D0 U3948 ( .A1(n7130), .A2(prog_data[3]), .B1(\mem[52][3] ), .B2(n7129), 
        .Z(n3824) );
  OA22D0 U3949 ( .A1(n7130), .A2(prog_data[2]), .B1(\mem[52][2] ), .B2(n7129), 
        .Z(n3823) );
  OA22D0 U3950 ( .A1(n7130), .A2(prog_data[1]), .B1(\mem[52][1] ), .B2(n7129), 
        .Z(n3822) );
  OA22D0 U3951 ( .A1(n7130), .A2(prog_data[0]), .B1(\mem[52][0] ), .B2(n7129), 
        .Z(n3821) );
  NR2D0 U3952 ( .A1(n7543), .A2(n7151), .ZN(n7131) );
  INVD0 U3953 ( .I(n7131), .ZN(n7132) );
  OA22D0 U3954 ( .A1(n7132), .A2(prog_data[15]), .B1(\mem[53][15] ), .B2(n7131), .Z(n3820) );
  OA22D0 U3955 ( .A1(n7132), .A2(prog_data[14]), .B1(\mem[53][14] ), .B2(n7131), .Z(n3819) );
  OA22D0 U3956 ( .A1(n7132), .A2(prog_data[13]), .B1(\mem[53][13] ), .B2(n7131), .Z(n3818) );
  OA22D0 U3957 ( .A1(n7132), .A2(prog_data[12]), .B1(\mem[53][12] ), .B2(n7131), .Z(n3817) );
  OA22D0 U3958 ( .A1(n7132), .A2(prog_data[11]), .B1(\mem[53][11] ), .B2(n7131), .Z(n3816) );
  OA22D0 U3959 ( .A1(n7132), .A2(prog_data[10]), .B1(\mem[53][10] ), .B2(n7131), .Z(n3815) );
  OA22D0 U3960 ( .A1(n7132), .A2(prog_data[9]), .B1(\mem[53][9] ), .B2(n7131), 
        .Z(n3814) );
  OA22D0 U3961 ( .A1(n7132), .A2(prog_data[8]), .B1(\mem[53][8] ), .B2(n7131), 
        .Z(n3813) );
  OA22D0 U3962 ( .A1(n7132), .A2(prog_data[7]), .B1(\mem[53][7] ), .B2(n7131), 
        .Z(n3812) );
  OA22D0 U3963 ( .A1(n7132), .A2(prog_data[6]), .B1(\mem[53][6] ), .B2(n7131), 
        .Z(n3811) );
  OA22D0 U3964 ( .A1(n7132), .A2(prog_data[5]), .B1(\mem[53][5] ), .B2(n7131), 
        .Z(n3810) );
  OA22D0 U3965 ( .A1(n7132), .A2(prog_data[4]), .B1(\mem[53][4] ), .B2(n7131), 
        .Z(n3809) );
  OA22D0 U3966 ( .A1(n7132), .A2(prog_data[3]), .B1(\mem[53][3] ), .B2(n7131), 
        .Z(n3808) );
  OA22D0 U3967 ( .A1(n7132), .A2(prog_data[2]), .B1(\mem[53][2] ), .B2(n7131), 
        .Z(n3807) );
  OA22D0 U3968 ( .A1(n7132), .A2(prog_data[1]), .B1(\mem[53][1] ), .B2(n7131), 
        .Z(n3806) );
  OA22D0 U3969 ( .A1(n7132), .A2(prog_data[0]), .B1(\mem[53][0] ), .B2(n7131), 
        .Z(n3805) );
  NR2D0 U3970 ( .A1(n7546), .A2(n7151), .ZN(n7133) );
  OA22D0 U3971 ( .A1(n7134), .A2(prog_data[15]), .B1(\mem[54][15] ), .B2(n7133), .Z(n3804) );
  OA22D0 U3972 ( .A1(n7134), .A2(prog_data[14]), .B1(\mem[54][14] ), .B2(n7133), .Z(n3803) );
  OA22D0 U3973 ( .A1(n7134), .A2(prog_data[13]), .B1(\mem[54][13] ), .B2(n7133), .Z(n3802) );
  OA22D0 U3974 ( .A1(n7134), .A2(prog_data[12]), .B1(\mem[54][12] ), .B2(n7133), .Z(n3801) );
  OA22D0 U3975 ( .A1(n7134), .A2(prog_data[11]), .B1(\mem[54][11] ), .B2(n7133), .Z(n3800) );
  OA22D0 U3976 ( .A1(n7134), .A2(prog_data[10]), .B1(\mem[54][10] ), .B2(n7133), .Z(n3799) );
  OA22D0 U3977 ( .A1(n7134), .A2(prog_data[9]), .B1(\mem[54][9] ), .B2(n7133), 
        .Z(n3798) );
  OA22D0 U3978 ( .A1(n7134), .A2(prog_data[8]), .B1(\mem[54][8] ), .B2(n7133), 
        .Z(n3797) );
  OA22D0 U3979 ( .A1(n7134), .A2(prog_data[7]), .B1(\mem[54][7] ), .B2(n7133), 
        .Z(n3796) );
  OA22D0 U3980 ( .A1(n7134), .A2(prog_data[6]), .B1(\mem[54][6] ), .B2(n7133), 
        .Z(n3795) );
  OA22D0 U3981 ( .A1(n7134), .A2(prog_data[5]), .B1(\mem[54][5] ), .B2(n7133), 
        .Z(n3794) );
  OA22D0 U3982 ( .A1(n7134), .A2(prog_data[4]), .B1(\mem[54][4] ), .B2(n7133), 
        .Z(n3793) );
  OA22D0 U3983 ( .A1(n7134), .A2(prog_data[3]), .B1(\mem[54][3] ), .B2(n7133), 
        .Z(n3792) );
  OA22D0 U3984 ( .A1(n7134), .A2(prog_data[2]), .B1(\mem[54][2] ), .B2(n7133), 
        .Z(n3791) );
  OA22D0 U3985 ( .A1(n7134), .A2(prog_data[1]), .B1(\mem[54][1] ), .B2(n7133), 
        .Z(n3790) );
  OA22D0 U3986 ( .A1(n7134), .A2(prog_data[0]), .B1(\mem[54][0] ), .B2(n7133), 
        .Z(n3789) );
  NR2D0 U3987 ( .A1(n7549), .A2(n7151), .ZN(n7135) );
  INVD0 U3988 ( .I(n7135), .ZN(n7136) );
  OA22D0 U3989 ( .A1(n7136), .A2(prog_data[15]), .B1(\mem[55][15] ), .B2(n7135), .Z(n3788) );
  OA22D0 U3990 ( .A1(n7136), .A2(prog_data[14]), .B1(\mem[55][14] ), .B2(n7135), .Z(n3787) );
  OA22D0 U3991 ( .A1(n7136), .A2(prog_data[13]), .B1(\mem[55][13] ), .B2(n7135), .Z(n3786) );
  OA22D0 U3992 ( .A1(n7136), .A2(prog_data[12]), .B1(\mem[55][12] ), .B2(n7135), .Z(n3785) );
  OA22D0 U3993 ( .A1(n7136), .A2(prog_data[11]), .B1(\mem[55][11] ), .B2(n7135), .Z(n3784) );
  OA22D0 U3994 ( .A1(n7136), .A2(prog_data[10]), .B1(\mem[55][10] ), .B2(n7135), .Z(n3783) );
  OA22D0 U3995 ( .A1(n7136), .A2(prog_data[9]), .B1(\mem[55][9] ), .B2(n7135), 
        .Z(n3782) );
  OA22D0 U3996 ( .A1(n7136), .A2(prog_data[8]), .B1(\mem[55][8] ), .B2(n7135), 
        .Z(n3781) );
  OA22D0 U3997 ( .A1(n7136), .A2(prog_data[7]), .B1(\mem[55][7] ), .B2(n7135), 
        .Z(n3780) );
  OA22D0 U3998 ( .A1(n7136), .A2(prog_data[6]), .B1(\mem[55][6] ), .B2(n7135), 
        .Z(n3779) );
  OA22D0 U3999 ( .A1(n7136), .A2(prog_data[5]), .B1(\mem[55][5] ), .B2(n7135), 
        .Z(n3778) );
  OA22D0 U4000 ( .A1(n7136), .A2(prog_data[4]), .B1(\mem[55][4] ), .B2(n7135), 
        .Z(n3777) );
  OA22D0 U4001 ( .A1(n7136), .A2(prog_data[3]), .B1(\mem[55][3] ), .B2(n7135), 
        .Z(n3776) );
  OA22D0 U4002 ( .A1(n7136), .A2(prog_data[2]), .B1(\mem[55][2] ), .B2(n7135), 
        .Z(n3775) );
  OA22D0 U4003 ( .A1(n7136), .A2(prog_data[1]), .B1(\mem[55][1] ), .B2(n7135), 
        .Z(n3774) );
  OA22D0 U4004 ( .A1(n7136), .A2(prog_data[0]), .B1(\mem[55][0] ), .B2(n7135), 
        .Z(n3773) );
  NR2D0 U4005 ( .A1(n7552), .A2(n7151), .ZN(n7137) );
  INVD0 U4006 ( .I(n7137), .ZN(n7138) );
  OA22D0 U4007 ( .A1(n7138), .A2(prog_data[15]), .B1(\mem[56][15] ), .B2(n7137), .Z(n3772) );
  OA22D0 U4008 ( .A1(n7138), .A2(prog_data[14]), .B1(\mem[56][14] ), .B2(n7137), .Z(n3771) );
  OA22D0 U4009 ( .A1(n7138), .A2(prog_data[13]), .B1(\mem[56][13] ), .B2(n7137), .Z(n3770) );
  OA22D0 U4010 ( .A1(n7138), .A2(prog_data[12]), .B1(\mem[56][12] ), .B2(n7137), .Z(n3769) );
  OA22D0 U4011 ( .A1(n7138), .A2(prog_data[11]), .B1(\mem[56][11] ), .B2(n7137), .Z(n3768) );
  OA22D0 U4012 ( .A1(n7138), .A2(prog_data[10]), .B1(\mem[56][10] ), .B2(n7137), .Z(n3767) );
  OA22D0 U4013 ( .A1(n7138), .A2(prog_data[9]), .B1(\mem[56][9] ), .B2(n7137), 
        .Z(n3766) );
  OA22D0 U4014 ( .A1(n7138), .A2(prog_data[8]), .B1(\mem[56][8] ), .B2(n7137), 
        .Z(n3765) );
  OA22D0 U4015 ( .A1(n7138), .A2(prog_data[7]), .B1(\mem[56][7] ), .B2(n7137), 
        .Z(n3764) );
  OA22D0 U4016 ( .A1(n7138), .A2(prog_data[6]), .B1(\mem[56][6] ), .B2(n7137), 
        .Z(n3763) );
  OA22D0 U4017 ( .A1(n7138), .A2(prog_data[5]), .B1(\mem[56][5] ), .B2(n7137), 
        .Z(n3762) );
  OA22D0 U4018 ( .A1(n7138), .A2(prog_data[4]), .B1(\mem[56][4] ), .B2(n7137), 
        .Z(n3761) );
  OA22D0 U4019 ( .A1(n7138), .A2(prog_data[3]), .B1(\mem[56][3] ), .B2(n7137), 
        .Z(n3760) );
  OA22D0 U4020 ( .A1(n7138), .A2(prog_data[2]), .B1(\mem[56][2] ), .B2(n7137), 
        .Z(n3759) );
  OA22D0 U4021 ( .A1(n7138), .A2(prog_data[1]), .B1(\mem[56][1] ), .B2(n7137), 
        .Z(n3758) );
  OA22D0 U4022 ( .A1(n7138), .A2(prog_data[0]), .B1(\mem[56][0] ), .B2(n7137), 
        .Z(n3757) );
  NR2D0 U4023 ( .A1(n7555), .A2(n7151), .ZN(n7139) );
  INVD0 U4024 ( .I(n7139), .ZN(n7140) );
  OA22D0 U4025 ( .A1(n7140), .A2(prog_data[15]), .B1(\mem[57][15] ), .B2(n7139), .Z(n3756) );
  OA22D0 U4026 ( .A1(n7140), .A2(prog_data[14]), .B1(\mem[57][14] ), .B2(n7139), .Z(n3755) );
  OA22D0 U4027 ( .A1(n7140), .A2(prog_data[13]), .B1(\mem[57][13] ), .B2(n7139), .Z(n3754) );
  OA22D0 U4028 ( .A1(n7140), .A2(prog_data[12]), .B1(\mem[57][12] ), .B2(n7139), .Z(n3753) );
  OA22D0 U4029 ( .A1(n7140), .A2(prog_data[11]), .B1(\mem[57][11] ), .B2(n7139), .Z(n3752) );
  OA22D0 U4030 ( .A1(n7140), .A2(prog_data[10]), .B1(\mem[57][10] ), .B2(n7139), .Z(n3751) );
  OA22D0 U4031 ( .A1(n7140), .A2(prog_data[9]), .B1(\mem[57][9] ), .B2(n7139), 
        .Z(n3750) );
  OA22D0 U4032 ( .A1(n7140), .A2(prog_data[8]), .B1(\mem[57][8] ), .B2(n7139), 
        .Z(n3749) );
  OA22D0 U4033 ( .A1(n7140), .A2(prog_data[7]), .B1(\mem[57][7] ), .B2(n7139), 
        .Z(n3748) );
  OA22D0 U4034 ( .A1(n7140), .A2(prog_data[6]), .B1(\mem[57][6] ), .B2(n7139), 
        .Z(n3747) );
  OA22D0 U4035 ( .A1(n7140), .A2(prog_data[5]), .B1(\mem[57][5] ), .B2(n7139), 
        .Z(n3746) );
  OA22D0 U4036 ( .A1(n7140), .A2(prog_data[4]), .B1(\mem[57][4] ), .B2(n7139), 
        .Z(n3745) );
  OA22D0 U4037 ( .A1(n7140), .A2(prog_data[3]), .B1(\mem[57][3] ), .B2(n7139), 
        .Z(n3744) );
  OA22D0 U4038 ( .A1(n7140), .A2(prog_data[2]), .B1(\mem[57][2] ), .B2(n7139), 
        .Z(n3743) );
  OA22D0 U4039 ( .A1(n7140), .A2(prog_data[1]), .B1(\mem[57][1] ), .B2(n7139), 
        .Z(n3742) );
  OA22D0 U4040 ( .A1(n7140), .A2(prog_data[0]), .B1(\mem[57][0] ), .B2(n7139), 
        .Z(n3741) );
  NR2D0 U4041 ( .A1(n7558), .A2(n7151), .ZN(n7141) );
  INVD0 U4042 ( .I(n7141), .ZN(n7142) );
  OA22D0 U4043 ( .A1(n7142), .A2(prog_data[15]), .B1(\mem[58][15] ), .B2(n7141), .Z(n3740) );
  OA22D0 U4044 ( .A1(n7142), .A2(prog_data[14]), .B1(\mem[58][14] ), .B2(n7141), .Z(n3739) );
  OA22D0 U4045 ( .A1(n7142), .A2(prog_data[13]), .B1(\mem[58][13] ), .B2(n7141), .Z(n3738) );
  OA22D0 U4046 ( .A1(n7142), .A2(prog_data[12]), .B1(\mem[58][12] ), .B2(n7141), .Z(n3737) );
  OA22D0 U4047 ( .A1(n7142), .A2(prog_data[11]), .B1(\mem[58][11] ), .B2(n7141), .Z(n3736) );
  OA22D0 U4048 ( .A1(n7142), .A2(prog_data[10]), .B1(\mem[58][10] ), .B2(n7141), .Z(n3735) );
  OA22D0 U4049 ( .A1(n7142), .A2(prog_data[9]), .B1(\mem[58][9] ), .B2(n7141), 
        .Z(n3734) );
  OA22D0 U4050 ( .A1(n7142), .A2(prog_data[8]), .B1(\mem[58][8] ), .B2(n7141), 
        .Z(n3733) );
  OA22D0 U4051 ( .A1(n7142), .A2(prog_data[7]), .B1(\mem[58][7] ), .B2(n7141), 
        .Z(n3732) );
  OA22D0 U4052 ( .A1(n7142), .A2(prog_data[6]), .B1(\mem[58][6] ), .B2(n7141), 
        .Z(n3731) );
  OA22D0 U4053 ( .A1(n7142), .A2(prog_data[5]), .B1(\mem[58][5] ), .B2(n7141), 
        .Z(n3730) );
  OA22D0 U4054 ( .A1(n7142), .A2(prog_data[4]), .B1(\mem[58][4] ), .B2(n7141), 
        .Z(n3729) );
  OA22D0 U4055 ( .A1(n7142), .A2(prog_data[3]), .B1(\mem[58][3] ), .B2(n7141), 
        .Z(n3728) );
  OA22D0 U4056 ( .A1(n7142), .A2(prog_data[2]), .B1(\mem[58][2] ), .B2(n7141), 
        .Z(n3727) );
  OA22D0 U4057 ( .A1(n7142), .A2(prog_data[1]), .B1(\mem[58][1] ), .B2(n7141), 
        .Z(n3726) );
  OA22D0 U4058 ( .A1(n7142), .A2(prog_data[0]), .B1(\mem[58][0] ), .B2(n7141), 
        .Z(n3725) );
  NR2D0 U4059 ( .A1(n7561), .A2(n7151), .ZN(n7143) );
  INVD0 U4060 ( .I(n7143), .ZN(n7144) );
  OA22D0 U4061 ( .A1(n7144), .A2(prog_data[15]), .B1(\mem[59][15] ), .B2(n7143), .Z(n3724) );
  OA22D0 U4062 ( .A1(n7144), .A2(prog_data[14]), .B1(\mem[59][14] ), .B2(n7143), .Z(n3723) );
  OA22D0 U4063 ( .A1(n7144), .A2(prog_data[13]), .B1(\mem[59][13] ), .B2(n7143), .Z(n3722) );
  OA22D0 U4064 ( .A1(n7144), .A2(prog_data[12]), .B1(\mem[59][12] ), .B2(n7143), .Z(n3721) );
  OA22D0 U4065 ( .A1(n7144), .A2(prog_data[11]), .B1(\mem[59][11] ), .B2(n7143), .Z(n3720) );
  OA22D0 U4066 ( .A1(n7144), .A2(prog_data[10]), .B1(\mem[59][10] ), .B2(n7143), .Z(n3719) );
  OA22D0 U4067 ( .A1(n7144), .A2(prog_data[9]), .B1(\mem[59][9] ), .B2(n7143), 
        .Z(n3718) );
  OA22D0 U4068 ( .A1(n7144), .A2(prog_data[8]), .B1(\mem[59][8] ), .B2(n7143), 
        .Z(n3717) );
  OA22D0 U4069 ( .A1(n7144), .A2(prog_data[7]), .B1(\mem[59][7] ), .B2(n7143), 
        .Z(n3716) );
  OA22D0 U4070 ( .A1(n7144), .A2(prog_data[6]), .B1(\mem[59][6] ), .B2(n7143), 
        .Z(n3715) );
  OA22D0 U4071 ( .A1(n7144), .A2(prog_data[5]), .B1(\mem[59][5] ), .B2(n7143), 
        .Z(n3714) );
  OA22D0 U4072 ( .A1(n7144), .A2(prog_data[4]), .B1(\mem[59][4] ), .B2(n7143), 
        .Z(n3713) );
  OA22D0 U4073 ( .A1(n7144), .A2(prog_data[3]), .B1(\mem[59][3] ), .B2(n7143), 
        .Z(n3712) );
  OA22D0 U4074 ( .A1(n7144), .A2(prog_data[2]), .B1(\mem[59][2] ), .B2(n7143), 
        .Z(n3711) );
  OA22D0 U4075 ( .A1(n7144), .A2(prog_data[1]), .B1(\mem[59][1] ), .B2(n7143), 
        .Z(n3710) );
  OA22D0 U4076 ( .A1(n7144), .A2(prog_data[0]), .B1(\mem[59][0] ), .B2(n7143), 
        .Z(n3709) );
  NR2D0 U4077 ( .A1(n7564), .A2(n7151), .ZN(n7145) );
  INVD0 U4078 ( .I(n7145), .ZN(n7146) );
  OA22D0 U4079 ( .A1(n7146), .A2(prog_data[15]), .B1(\mem[60][15] ), .B2(n7145), .Z(n3708) );
  OA22D0 U4080 ( .A1(n7146), .A2(prog_data[14]), .B1(\mem[60][14] ), .B2(n7145), .Z(n3707) );
  OA22D0 U4081 ( .A1(n7146), .A2(prog_data[13]), .B1(\mem[60][13] ), .B2(n7145), .Z(n3706) );
  OA22D0 U4082 ( .A1(n7146), .A2(prog_data[12]), .B1(\mem[60][12] ), .B2(n7145), .Z(n3705) );
  OA22D0 U4083 ( .A1(n7146), .A2(prog_data[11]), .B1(\mem[60][11] ), .B2(n7145), .Z(n3704) );
  OA22D0 U4084 ( .A1(n7146), .A2(prog_data[10]), .B1(\mem[60][10] ), .B2(n7145), .Z(n3703) );
  OA22D0 U4085 ( .A1(n7146), .A2(prog_data[9]), .B1(\mem[60][9] ), .B2(n7145), 
        .Z(n3702) );
  OA22D0 U4086 ( .A1(n7146), .A2(prog_data[8]), .B1(\mem[60][8] ), .B2(n7145), 
        .Z(n3701) );
  OA22D0 U4087 ( .A1(n7146), .A2(prog_data[7]), .B1(\mem[60][7] ), .B2(n7145), 
        .Z(n3700) );
  OA22D0 U4088 ( .A1(n7146), .A2(prog_data[6]), .B1(\mem[60][6] ), .B2(n7145), 
        .Z(n3699) );
  OA22D0 U4089 ( .A1(n7146), .A2(prog_data[5]), .B1(\mem[60][5] ), .B2(n7145), 
        .Z(n3698) );
  OA22D0 U4090 ( .A1(n7146), .A2(prog_data[4]), .B1(\mem[60][4] ), .B2(n7145), 
        .Z(n3697) );
  OA22D0 U4091 ( .A1(n7146), .A2(prog_data[3]), .B1(\mem[60][3] ), .B2(n7145), 
        .Z(n3696) );
  OA22D0 U4092 ( .A1(n7146), .A2(prog_data[2]), .B1(\mem[60][2] ), .B2(n7145), 
        .Z(n3695) );
  OA22D0 U4093 ( .A1(n7146), .A2(prog_data[1]), .B1(\mem[60][1] ), .B2(n7145), 
        .Z(n3694) );
  OA22D0 U4094 ( .A1(n7146), .A2(prog_data[0]), .B1(\mem[60][0] ), .B2(n7145), 
        .Z(n3693) );
  INVD0 U4095 ( .I(n7147), .ZN(n7148) );
  OA22D0 U4096 ( .A1(n7148), .A2(prog_data[15]), .B1(\mem[61][15] ), .B2(n7147), .Z(n3692) );
  OA22D0 U4097 ( .A1(n7148), .A2(prog_data[14]), .B1(\mem[61][14] ), .B2(n7147), .Z(n3691) );
  OA22D0 U4098 ( .A1(n7148), .A2(prog_data[13]), .B1(\mem[61][13] ), .B2(n7147), .Z(n3690) );
  OA22D0 U4099 ( .A1(n7148), .A2(prog_data[12]), .B1(\mem[61][12] ), .B2(n7147), .Z(n3689) );
  OA22D0 U4100 ( .A1(n7148), .A2(prog_data[11]), .B1(\mem[61][11] ), .B2(n7147), .Z(n3688) );
  OA22D0 U4101 ( .A1(n7148), .A2(prog_data[10]), .B1(\mem[61][10] ), .B2(n7147), .Z(n3687) );
  OA22D0 U4102 ( .A1(n7148), .A2(prog_data[9]), .B1(\mem[61][9] ), .B2(n7147), 
        .Z(n3686) );
  OA22D0 U4103 ( .A1(n7148), .A2(prog_data[8]), .B1(\mem[61][8] ), .B2(n7147), 
        .Z(n3685) );
  OA22D0 U4104 ( .A1(n7148), .A2(prog_data[7]), .B1(\mem[61][7] ), .B2(n7147), 
        .Z(n3684) );
  OA22D0 U4105 ( .A1(n7148), .A2(prog_data[6]), .B1(\mem[61][6] ), .B2(n7147), 
        .Z(n3683) );
  OA22D0 U4106 ( .A1(n7148), .A2(prog_data[5]), .B1(\mem[61][5] ), .B2(n7147), 
        .Z(n3682) );
  OA22D0 U4107 ( .A1(n7148), .A2(prog_data[4]), .B1(\mem[61][4] ), .B2(n7147), 
        .Z(n3681) );
  OA22D0 U4108 ( .A1(n7148), .A2(prog_data[3]), .B1(\mem[61][3] ), .B2(n7147), 
        .Z(n3680) );
  OA22D0 U4109 ( .A1(n7148), .A2(prog_data[2]), .B1(\mem[61][2] ), .B2(n7147), 
        .Z(n3679) );
  OA22D0 U4110 ( .A1(n7148), .A2(prog_data[1]), .B1(\mem[61][1] ), .B2(n7147), 
        .Z(n3678) );
  OA22D0 U4111 ( .A1(n7148), .A2(prog_data[0]), .B1(\mem[61][0] ), .B2(n7147), 
        .Z(n3677) );
  NR2D0 U4112 ( .A1(n7570), .A2(n7151), .ZN(n7149) );
  INVD0 U4113 ( .I(n7149), .ZN(n7150) );
  OA22D0 U4114 ( .A1(n7150), .A2(prog_data[15]), .B1(\mem[62][15] ), .B2(n7149), .Z(n3676) );
  OA22D0 U4115 ( .A1(n7150), .A2(prog_data[14]), .B1(\mem[62][14] ), .B2(n7149), .Z(n3675) );
  OA22D0 U4116 ( .A1(n7150), .A2(prog_data[13]), .B1(\mem[62][13] ), .B2(n7149), .Z(n3674) );
  OA22D0 U4117 ( .A1(n7150), .A2(prog_data[12]), .B1(\mem[62][12] ), .B2(n7149), .Z(n3673) );
  OA22D0 U4118 ( .A1(n7150), .A2(prog_data[11]), .B1(\mem[62][11] ), .B2(n7149), .Z(n3672) );
  OA22D0 U4119 ( .A1(n7150), .A2(prog_data[10]), .B1(\mem[62][10] ), .B2(n7149), .Z(n3671) );
  OA22D0 U4120 ( .A1(n7150), .A2(prog_data[9]), .B1(\mem[62][9] ), .B2(n7149), 
        .Z(n3670) );
  OA22D0 U4121 ( .A1(n7150), .A2(prog_data[8]), .B1(\mem[62][8] ), .B2(n7149), 
        .Z(n3669) );
  OA22D0 U4122 ( .A1(n7150), .A2(prog_data[7]), .B1(\mem[62][7] ), .B2(n7149), 
        .Z(n3668) );
  OA22D0 U4123 ( .A1(n7150), .A2(prog_data[6]), .B1(\mem[62][6] ), .B2(n7149), 
        .Z(n3667) );
  OA22D0 U4124 ( .A1(n7150), .A2(prog_data[5]), .B1(\mem[62][5] ), .B2(n7149), 
        .Z(n3666) );
  OA22D0 U4125 ( .A1(n7150), .A2(prog_data[4]), .B1(\mem[62][4] ), .B2(n7149), 
        .Z(n3665) );
  OA22D0 U4126 ( .A1(n7150), .A2(prog_data[3]), .B1(\mem[62][3] ), .B2(n7149), 
        .Z(n3664) );
  OA22D0 U4127 ( .A1(n7150), .A2(prog_data[2]), .B1(\mem[62][2] ), .B2(n7149), 
        .Z(n3663) );
  OA22D0 U4128 ( .A1(n7150), .A2(prog_data[1]), .B1(\mem[62][1] ), .B2(n7149), 
        .Z(n3662) );
  OA22D0 U4129 ( .A1(n7150), .A2(prog_data[0]), .B1(\mem[62][0] ), .B2(n7149), 
        .Z(n3661) );
  NR2D0 U4130 ( .A1(n7574), .A2(n7151), .ZN(n7152) );
  INVD0 U4131 ( .I(n7152), .ZN(n7153) );
  OA22D0 U4132 ( .A1(n7153), .A2(prog_data[15]), .B1(\mem[63][15] ), .B2(n7152), .Z(n3660) );
  OA22D0 U4133 ( .A1(n7153), .A2(prog_data[14]), .B1(\mem[63][14] ), .B2(n7152), .Z(n3659) );
  OA22D0 U4134 ( .A1(n7153), .A2(prog_data[13]), .B1(\mem[63][13] ), .B2(n7152), .Z(n3658) );
  OA22D0 U4135 ( .A1(n7153), .A2(prog_data[12]), .B1(\mem[63][12] ), .B2(n7152), .Z(n3657) );
  OA22D0 U4136 ( .A1(n7153), .A2(prog_data[11]), .B1(\mem[63][11] ), .B2(n7152), .Z(n3656) );
  OA22D0 U4137 ( .A1(n7153), .A2(prog_data[10]), .B1(\mem[63][10] ), .B2(n7152), .Z(n3655) );
  OA22D0 U4138 ( .A1(n7153), .A2(prog_data[9]), .B1(\mem[63][9] ), .B2(n7152), 
        .Z(n3654) );
  OA22D0 U4139 ( .A1(n7153), .A2(prog_data[8]), .B1(\mem[63][8] ), .B2(n7152), 
        .Z(n3653) );
  OA22D0 U4140 ( .A1(n7153), .A2(prog_data[7]), .B1(\mem[63][7] ), .B2(n7152), 
        .Z(n3652) );
  OA22D0 U4141 ( .A1(n7153), .A2(prog_data[6]), .B1(\mem[63][6] ), .B2(n7152), 
        .Z(n3651) );
  OA22D0 U4142 ( .A1(n7153), .A2(prog_data[5]), .B1(\mem[63][5] ), .B2(n7152), 
        .Z(n3650) );
  OA22D0 U4143 ( .A1(n7153), .A2(prog_data[4]), .B1(\mem[63][4] ), .B2(n7152), 
        .Z(n3649) );
  OA22D0 U4144 ( .A1(n7153), .A2(prog_data[3]), .B1(\mem[63][3] ), .B2(n7152), 
        .Z(n3648) );
  OA22D0 U4145 ( .A1(n7153), .A2(prog_data[2]), .B1(\mem[63][2] ), .B2(n7152), 
        .Z(n3647) );
  OA22D0 U4146 ( .A1(n7153), .A2(prog_data[1]), .B1(\mem[63][1] ), .B2(n7152), 
        .Z(n3646) );
  OA22D0 U4147 ( .A1(n7153), .A2(prog_data[0]), .B1(\mem[63][0] ), .B2(n7152), 
        .Z(n3645) );
  ND3D0 U4148 ( .A1(prog_addr[6]), .A2(n7221), .A3(n7187), .ZN(n7184) );
  NR2D0 U4149 ( .A1(n7528), .A2(n7184), .ZN(n7154) );
  INVD0 U4150 ( .I(n7154), .ZN(n7155) );
  OA22D0 U4151 ( .A1(n7155), .A2(prog_data[15]), .B1(\mem[64][15] ), .B2(n7154), .Z(n3644) );
  OA22D0 U4152 ( .A1(n7155), .A2(prog_data[14]), .B1(\mem[64][14] ), .B2(n7154), .Z(n3643) );
  OA22D0 U4153 ( .A1(n7155), .A2(prog_data[13]), .B1(\mem[64][13] ), .B2(n7154), .Z(n3642) );
  OA22D0 U4154 ( .A1(n7155), .A2(prog_data[12]), .B1(\mem[64][12] ), .B2(n7154), .Z(n3641) );
  OA22D0 U4155 ( .A1(n7155), .A2(prog_data[11]), .B1(\mem[64][11] ), .B2(n7154), .Z(n3640) );
  OA22D0 U4156 ( .A1(n7155), .A2(prog_data[10]), .B1(\mem[64][10] ), .B2(n7154), .Z(n3639) );
  OA22D0 U4157 ( .A1(n7155), .A2(prog_data[9]), .B1(\mem[64][9] ), .B2(n7154), 
        .Z(n3638) );
  OA22D0 U4158 ( .A1(n7155), .A2(prog_data[8]), .B1(\mem[64][8] ), .B2(n7154), 
        .Z(n3637) );
  OA22D0 U4159 ( .A1(n7155), .A2(prog_data[7]), .B1(\mem[64][7] ), .B2(n7154), 
        .Z(n3636) );
  OA22D0 U4160 ( .A1(n7155), .A2(prog_data[6]), .B1(\mem[64][6] ), .B2(n7154), 
        .Z(n3635) );
  OA22D0 U4161 ( .A1(n7155), .A2(prog_data[5]), .B1(\mem[64][5] ), .B2(n7154), 
        .Z(n3634) );
  OA22D0 U4162 ( .A1(n7155), .A2(prog_data[4]), .B1(\mem[64][4] ), .B2(n7154), 
        .Z(n3633) );
  OA22D0 U4163 ( .A1(n7155), .A2(prog_data[3]), .B1(\mem[64][3] ), .B2(n7154), 
        .Z(n3632) );
  OA22D0 U4164 ( .A1(n7155), .A2(prog_data[2]), .B1(\mem[64][2] ), .B2(n7154), 
        .Z(n3631) );
  OA22D0 U4165 ( .A1(n7155), .A2(prog_data[1]), .B1(\mem[64][1] ), .B2(n7154), 
        .Z(n3630) );
  OA22D0 U4166 ( .A1(n7155), .A2(prog_data[0]), .B1(\mem[64][0] ), .B2(n7154), 
        .Z(n3629) );
  NR2D0 U4167 ( .A1(n7531), .A2(n7184), .ZN(n7156) );
  INVD0 U4168 ( .I(n7156), .ZN(n7157) );
  OA22D0 U4169 ( .A1(n7157), .A2(prog_data[15]), .B1(\mem[65][15] ), .B2(n7156), .Z(n3628) );
  OA22D0 U4170 ( .A1(n7157), .A2(prog_data[14]), .B1(\mem[65][14] ), .B2(n7156), .Z(n3627) );
  OA22D0 U4171 ( .A1(n7157), .A2(prog_data[13]), .B1(\mem[65][13] ), .B2(n7156), .Z(n3626) );
  OA22D0 U4172 ( .A1(n7157), .A2(prog_data[12]), .B1(\mem[65][12] ), .B2(n7156), .Z(n3625) );
  OA22D0 U4173 ( .A1(n7157), .A2(prog_data[11]), .B1(\mem[65][11] ), .B2(n7156), .Z(n3624) );
  OA22D0 U4174 ( .A1(n7157), .A2(prog_data[10]), .B1(\mem[65][10] ), .B2(n7156), .Z(n3623) );
  OA22D0 U4175 ( .A1(n7157), .A2(prog_data[9]), .B1(\mem[65][9] ), .B2(n7156), 
        .Z(n3622) );
  OA22D0 U4176 ( .A1(n7157), .A2(prog_data[8]), .B1(\mem[65][8] ), .B2(n7156), 
        .Z(n3621) );
  OA22D0 U4177 ( .A1(n7157), .A2(prog_data[7]), .B1(\mem[65][7] ), .B2(n7156), 
        .Z(n3620) );
  OA22D0 U4178 ( .A1(n7157), .A2(prog_data[6]), .B1(\mem[65][6] ), .B2(n7156), 
        .Z(n3619) );
  OA22D0 U4179 ( .A1(n7157), .A2(prog_data[5]), .B1(\mem[65][5] ), .B2(n7156), 
        .Z(n3618) );
  OA22D0 U4180 ( .A1(n7157), .A2(prog_data[4]), .B1(\mem[65][4] ), .B2(n7156), 
        .Z(n3617) );
  OA22D0 U4181 ( .A1(n7157), .A2(prog_data[3]), .B1(\mem[65][3] ), .B2(n7156), 
        .Z(n3616) );
  OA22D0 U4182 ( .A1(n7157), .A2(prog_data[2]), .B1(\mem[65][2] ), .B2(n7156), 
        .Z(n3615) );
  OA22D0 U4183 ( .A1(n7157), .A2(prog_data[1]), .B1(\mem[65][1] ), .B2(n7156), 
        .Z(n3614) );
  OA22D0 U4184 ( .A1(n7157), .A2(prog_data[0]), .B1(\mem[65][0] ), .B2(n7156), 
        .Z(n3613) );
  NR2D0 U4185 ( .A1(n7534), .A2(n7184), .ZN(n7158) );
  INVD0 U4186 ( .I(n7158), .ZN(n7159) );
  OA22D0 U4187 ( .A1(n7159), .A2(prog_data[15]), .B1(\mem[66][15] ), .B2(n7158), .Z(n3612) );
  OA22D0 U4188 ( .A1(n7159), .A2(prog_data[14]), .B1(\mem[66][14] ), .B2(n7158), .Z(n3611) );
  OA22D0 U4189 ( .A1(n7159), .A2(prog_data[13]), .B1(\mem[66][13] ), .B2(n7158), .Z(n3610) );
  OA22D0 U4190 ( .A1(n7159), .A2(prog_data[12]), .B1(\mem[66][12] ), .B2(n7158), .Z(n3609) );
  OA22D0 U4191 ( .A1(n7159), .A2(prog_data[11]), .B1(\mem[66][11] ), .B2(n7158), .Z(n3608) );
  OA22D0 U4192 ( .A1(n7159), .A2(prog_data[10]), .B1(\mem[66][10] ), .B2(n7158), .Z(n3607) );
  OA22D0 U4193 ( .A1(n7159), .A2(prog_data[9]), .B1(\mem[66][9] ), .B2(n7158), 
        .Z(n3606) );
  OA22D0 U4194 ( .A1(n7159), .A2(prog_data[8]), .B1(\mem[66][8] ), .B2(n7158), 
        .Z(n3605) );
  OA22D0 U4195 ( .A1(n7159), .A2(prog_data[7]), .B1(\mem[66][7] ), .B2(n7158), 
        .Z(n3604) );
  OA22D0 U4196 ( .A1(n7159), .A2(prog_data[6]), .B1(\mem[66][6] ), .B2(n7158), 
        .Z(n3603) );
  OA22D0 U4197 ( .A1(n7159), .A2(prog_data[5]), .B1(\mem[66][5] ), .B2(n7158), 
        .Z(n3602) );
  OA22D0 U4198 ( .A1(n7159), .A2(prog_data[4]), .B1(\mem[66][4] ), .B2(n7158), 
        .Z(n3601) );
  OA22D0 U4199 ( .A1(n7159), .A2(prog_data[3]), .B1(\mem[66][3] ), .B2(n7158), 
        .Z(n3600) );
  OA22D0 U4200 ( .A1(n7159), .A2(prog_data[2]), .B1(\mem[66][2] ), .B2(n7158), 
        .Z(n3599) );
  OA22D0 U4201 ( .A1(n7159), .A2(prog_data[1]), .B1(\mem[66][1] ), .B2(n7158), 
        .Z(n3598) );
  OA22D0 U4202 ( .A1(n7159), .A2(prog_data[0]), .B1(\mem[66][0] ), .B2(n7158), 
        .Z(n3597) );
  NR2D0 U4203 ( .A1(n7537), .A2(n7184), .ZN(n7160) );
  INVD0 U4204 ( .I(n7160), .ZN(n7161) );
  OA22D0 U4205 ( .A1(n7161), .A2(prog_data[15]), .B1(\mem[67][15] ), .B2(n7160), .Z(n3596) );
  OA22D0 U4206 ( .A1(n7161), .A2(prog_data[14]), .B1(\mem[67][14] ), .B2(n7160), .Z(n3595) );
  OA22D0 U4207 ( .A1(n7161), .A2(prog_data[13]), .B1(\mem[67][13] ), .B2(n7160), .Z(n3594) );
  OA22D0 U4208 ( .A1(n7161), .A2(prog_data[12]), .B1(\mem[67][12] ), .B2(n7160), .Z(n3593) );
  OA22D0 U4209 ( .A1(n7161), .A2(prog_data[11]), .B1(\mem[67][11] ), .B2(n7160), .Z(n3592) );
  OA22D0 U4210 ( .A1(n7161), .A2(prog_data[10]), .B1(\mem[67][10] ), .B2(n7160), .Z(n3591) );
  OA22D0 U4211 ( .A1(n7161), .A2(prog_data[9]), .B1(\mem[67][9] ), .B2(n7160), 
        .Z(n3590) );
  OA22D0 U4212 ( .A1(n7161), .A2(prog_data[8]), .B1(\mem[67][8] ), .B2(n7160), 
        .Z(n3589) );
  OA22D0 U4213 ( .A1(n7161), .A2(prog_data[7]), .B1(\mem[67][7] ), .B2(n7160), 
        .Z(n3588) );
  OA22D0 U4214 ( .A1(n7161), .A2(prog_data[6]), .B1(\mem[67][6] ), .B2(n7160), 
        .Z(n3587) );
  OA22D0 U4215 ( .A1(n7161), .A2(prog_data[5]), .B1(\mem[67][5] ), .B2(n7160), 
        .Z(n3586) );
  OA22D0 U4216 ( .A1(n7161), .A2(prog_data[4]), .B1(\mem[67][4] ), .B2(n7160), 
        .Z(n3585) );
  OA22D0 U4217 ( .A1(n7161), .A2(prog_data[3]), .B1(\mem[67][3] ), .B2(n7160), 
        .Z(n3584) );
  OA22D0 U4218 ( .A1(n7161), .A2(prog_data[2]), .B1(\mem[67][2] ), .B2(n7160), 
        .Z(n3583) );
  OA22D0 U4219 ( .A1(n7161), .A2(prog_data[1]), .B1(\mem[67][1] ), .B2(n7160), 
        .Z(n3582) );
  OA22D0 U4220 ( .A1(n7161), .A2(prog_data[0]), .B1(\mem[67][0] ), .B2(n7160), 
        .Z(n3581) );
  NR2D0 U4221 ( .A1(n7540), .A2(n7184), .ZN(n7162) );
  INVD0 U4222 ( .I(n7162), .ZN(n7163) );
  OA22D0 U4223 ( .A1(n7163), .A2(prog_data[15]), .B1(\mem[68][15] ), .B2(n7162), .Z(n3580) );
  OA22D0 U4224 ( .A1(n7163), .A2(prog_data[14]), .B1(\mem[68][14] ), .B2(n7162), .Z(n3579) );
  OA22D0 U4225 ( .A1(n7163), .A2(prog_data[13]), .B1(\mem[68][13] ), .B2(n7162), .Z(n3578) );
  OA22D0 U4226 ( .A1(n7163), .A2(prog_data[12]), .B1(\mem[68][12] ), .B2(n7162), .Z(n3577) );
  OA22D0 U4227 ( .A1(n7163), .A2(prog_data[11]), .B1(\mem[68][11] ), .B2(n7162), .Z(n3576) );
  OA22D0 U4228 ( .A1(n7163), .A2(prog_data[10]), .B1(\mem[68][10] ), .B2(n7162), .Z(n3575) );
  OA22D0 U4229 ( .A1(n7163), .A2(prog_data[9]), .B1(\mem[68][9] ), .B2(n7162), 
        .Z(n3574) );
  OA22D0 U4230 ( .A1(n7163), .A2(prog_data[8]), .B1(\mem[68][8] ), .B2(n7162), 
        .Z(n3573) );
  OA22D0 U4231 ( .A1(n7163), .A2(prog_data[7]), .B1(\mem[68][7] ), .B2(n7162), 
        .Z(n3572) );
  OA22D0 U4232 ( .A1(n7163), .A2(prog_data[6]), .B1(\mem[68][6] ), .B2(n7162), 
        .Z(n3571) );
  OA22D0 U4233 ( .A1(n7163), .A2(prog_data[5]), .B1(\mem[68][5] ), .B2(n7162), 
        .Z(n3570) );
  OA22D0 U4234 ( .A1(n7163), .A2(prog_data[4]), .B1(\mem[68][4] ), .B2(n7162), 
        .Z(n3569) );
  OA22D0 U4235 ( .A1(n7163), .A2(prog_data[3]), .B1(\mem[68][3] ), .B2(n7162), 
        .Z(n3568) );
  OA22D0 U4236 ( .A1(n7163), .A2(prog_data[2]), .B1(\mem[68][2] ), .B2(n7162), 
        .Z(n3567) );
  OA22D0 U4237 ( .A1(n7163), .A2(prog_data[1]), .B1(\mem[68][1] ), .B2(n7162), 
        .Z(n3566) );
  OA22D0 U4238 ( .A1(n7163), .A2(prog_data[0]), .B1(\mem[68][0] ), .B2(n7162), 
        .Z(n3565) );
  NR2D0 U4239 ( .A1(n7543), .A2(n7184), .ZN(n7164) );
  OA22D0 U4240 ( .A1(n7165), .A2(prog_data[15]), .B1(\mem[69][15] ), .B2(n7164), .Z(n3564) );
  OA22D0 U4241 ( .A1(n7165), .A2(prog_data[14]), .B1(\mem[69][14] ), .B2(n7164), .Z(n3563) );
  OA22D0 U4242 ( .A1(n7165), .A2(prog_data[13]), .B1(\mem[69][13] ), .B2(n7164), .Z(n3562) );
  OA22D0 U4243 ( .A1(n7165), .A2(prog_data[12]), .B1(\mem[69][12] ), .B2(n7164), .Z(n3561) );
  OA22D0 U4244 ( .A1(n7165), .A2(prog_data[11]), .B1(\mem[69][11] ), .B2(n7164), .Z(n3560) );
  OA22D0 U4245 ( .A1(n7165), .A2(prog_data[10]), .B1(\mem[69][10] ), .B2(n7164), .Z(n3559) );
  OA22D0 U4246 ( .A1(n7165), .A2(prog_data[9]), .B1(\mem[69][9] ), .B2(n7164), 
        .Z(n3558) );
  OA22D0 U4247 ( .A1(n7165), .A2(prog_data[8]), .B1(\mem[69][8] ), .B2(n7164), 
        .Z(n3557) );
  OA22D0 U4248 ( .A1(n7165), .A2(prog_data[7]), .B1(\mem[69][7] ), .B2(n7164), 
        .Z(n3556) );
  OA22D0 U4249 ( .A1(n7165), .A2(prog_data[6]), .B1(\mem[69][6] ), .B2(n7164), 
        .Z(n3555) );
  OA22D0 U4250 ( .A1(n7165), .A2(prog_data[5]), .B1(\mem[69][5] ), .B2(n7164), 
        .Z(n3554) );
  OA22D0 U4251 ( .A1(n7165), .A2(prog_data[4]), .B1(\mem[69][4] ), .B2(n7164), 
        .Z(n3553) );
  OA22D0 U4252 ( .A1(n7165), .A2(prog_data[3]), .B1(\mem[69][3] ), .B2(n7164), 
        .Z(n3552) );
  OA22D0 U4253 ( .A1(n7165), .A2(prog_data[2]), .B1(\mem[69][2] ), .B2(n7164), 
        .Z(n3551) );
  OA22D0 U4254 ( .A1(n7165), .A2(prog_data[1]), .B1(\mem[69][1] ), .B2(n7164), 
        .Z(n3550) );
  OA22D0 U4255 ( .A1(n7165), .A2(prog_data[0]), .B1(\mem[69][0] ), .B2(n7164), 
        .Z(n3549) );
  NR2D0 U4256 ( .A1(n7546), .A2(n7184), .ZN(n7166) );
  INVD0 U4257 ( .I(n7166), .ZN(n7167) );
  OA22D0 U4258 ( .A1(n7167), .A2(prog_data[15]), .B1(\mem[70][15] ), .B2(n7166), .Z(n3548) );
  OA22D0 U4259 ( .A1(n7167), .A2(prog_data[14]), .B1(\mem[70][14] ), .B2(n7166), .Z(n3547) );
  OA22D0 U4260 ( .A1(n7167), .A2(prog_data[13]), .B1(\mem[70][13] ), .B2(n7166), .Z(n3546) );
  OA22D0 U4261 ( .A1(n7167), .A2(prog_data[12]), .B1(\mem[70][12] ), .B2(n7166), .Z(n3545) );
  OA22D0 U4262 ( .A1(n7167), .A2(prog_data[11]), .B1(\mem[70][11] ), .B2(n7166), .Z(n3544) );
  OA22D0 U4263 ( .A1(n7167), .A2(prog_data[10]), .B1(\mem[70][10] ), .B2(n7166), .Z(n3543) );
  OA22D0 U4264 ( .A1(n7167), .A2(prog_data[9]), .B1(\mem[70][9] ), .B2(n7166), 
        .Z(n3542) );
  OA22D0 U4265 ( .A1(n7167), .A2(prog_data[8]), .B1(\mem[70][8] ), .B2(n7166), 
        .Z(n3541) );
  OA22D0 U4266 ( .A1(n7167), .A2(prog_data[7]), .B1(\mem[70][7] ), .B2(n7166), 
        .Z(n3540) );
  OA22D0 U4267 ( .A1(n7167), .A2(prog_data[6]), .B1(\mem[70][6] ), .B2(n7166), 
        .Z(n3539) );
  OA22D0 U4268 ( .A1(n7167), .A2(prog_data[5]), .B1(\mem[70][5] ), .B2(n7166), 
        .Z(n3538) );
  OA22D0 U4269 ( .A1(n7167), .A2(prog_data[4]), .B1(\mem[70][4] ), .B2(n7166), 
        .Z(n3537) );
  OA22D0 U4270 ( .A1(n7167), .A2(prog_data[3]), .B1(\mem[70][3] ), .B2(n7166), 
        .Z(n3536) );
  OA22D0 U4271 ( .A1(n7167), .A2(prog_data[2]), .B1(\mem[70][2] ), .B2(n7166), 
        .Z(n3535) );
  OA22D0 U4272 ( .A1(n7167), .A2(prog_data[1]), .B1(\mem[70][1] ), .B2(n7166), 
        .Z(n3534) );
  OA22D0 U4273 ( .A1(n7167), .A2(prog_data[0]), .B1(\mem[70][0] ), .B2(n7166), 
        .Z(n3533) );
  NR2D0 U4274 ( .A1(n7549), .A2(n7184), .ZN(n7168) );
  INVD0 U4275 ( .I(n7168), .ZN(n7169) );
  OA22D0 U4276 ( .A1(n7169), .A2(prog_data[15]), .B1(\mem[71][15] ), .B2(n7168), .Z(n3532) );
  OA22D0 U4277 ( .A1(n7169), .A2(prog_data[14]), .B1(\mem[71][14] ), .B2(n7168), .Z(n3531) );
  OA22D0 U4278 ( .A1(n7169), .A2(prog_data[13]), .B1(\mem[71][13] ), .B2(n7168), .Z(n3530) );
  OA22D0 U4279 ( .A1(n7169), .A2(prog_data[12]), .B1(\mem[71][12] ), .B2(n7168), .Z(n3529) );
  OA22D0 U4280 ( .A1(n7169), .A2(prog_data[11]), .B1(\mem[71][11] ), .B2(n7168), .Z(n3528) );
  OA22D0 U4281 ( .A1(n7169), .A2(prog_data[10]), .B1(\mem[71][10] ), .B2(n7168), .Z(n3527) );
  OA22D0 U4282 ( .A1(n7169), .A2(prog_data[9]), .B1(\mem[71][9] ), .B2(n7168), 
        .Z(n3526) );
  OA22D0 U4283 ( .A1(n7169), .A2(prog_data[8]), .B1(\mem[71][8] ), .B2(n7168), 
        .Z(n3525) );
  OA22D0 U4284 ( .A1(n7169), .A2(prog_data[7]), .B1(\mem[71][7] ), .B2(n7168), 
        .Z(n3524) );
  OA22D0 U4285 ( .A1(n7169), .A2(prog_data[6]), .B1(\mem[71][6] ), .B2(n7168), 
        .Z(n3523) );
  OA22D0 U4286 ( .A1(n7169), .A2(prog_data[5]), .B1(\mem[71][5] ), .B2(n7168), 
        .Z(n3522) );
  OA22D0 U4287 ( .A1(n7169), .A2(prog_data[4]), .B1(\mem[71][4] ), .B2(n7168), 
        .Z(n3521) );
  OA22D0 U4288 ( .A1(n7169), .A2(prog_data[3]), .B1(\mem[71][3] ), .B2(n7168), 
        .Z(n3520) );
  OA22D0 U4289 ( .A1(n7169), .A2(prog_data[2]), .B1(\mem[71][2] ), .B2(n7168), 
        .Z(n3519) );
  OA22D0 U4290 ( .A1(n7169), .A2(prog_data[1]), .B1(\mem[71][1] ), .B2(n7168), 
        .Z(n3518) );
  OA22D0 U4291 ( .A1(n7169), .A2(prog_data[0]), .B1(\mem[71][0] ), .B2(n7168), 
        .Z(n3517) );
  NR2D0 U4292 ( .A1(n7552), .A2(n7184), .ZN(n7170) );
  INVD0 U4293 ( .I(n7170), .ZN(n7171) );
  OA22D0 U4294 ( .A1(n7171), .A2(prog_data[15]), .B1(\mem[72][15] ), .B2(n7170), .Z(n3516) );
  OA22D0 U4295 ( .A1(n7171), .A2(prog_data[14]), .B1(\mem[72][14] ), .B2(n7170), .Z(n3515) );
  OA22D0 U4296 ( .A1(n7171), .A2(prog_data[13]), .B1(\mem[72][13] ), .B2(n7170), .Z(n3514) );
  OA22D0 U4297 ( .A1(n7171), .A2(prog_data[12]), .B1(\mem[72][12] ), .B2(n7170), .Z(n3513) );
  OA22D0 U4298 ( .A1(n7171), .A2(prog_data[11]), .B1(\mem[72][11] ), .B2(n7170), .Z(n3512) );
  OA22D0 U4299 ( .A1(n7171), .A2(prog_data[10]), .B1(\mem[72][10] ), .B2(n7170), .Z(n3511) );
  OA22D0 U4300 ( .A1(n7171), .A2(prog_data[9]), .B1(\mem[72][9] ), .B2(n7170), 
        .Z(n3510) );
  OA22D0 U4301 ( .A1(n7171), .A2(prog_data[8]), .B1(\mem[72][8] ), .B2(n7170), 
        .Z(n3509) );
  OA22D0 U4302 ( .A1(n7171), .A2(prog_data[7]), .B1(\mem[72][7] ), .B2(n7170), 
        .Z(n3508) );
  OA22D0 U4303 ( .A1(n7171), .A2(prog_data[6]), .B1(\mem[72][6] ), .B2(n7170), 
        .Z(n3507) );
  OA22D0 U4304 ( .A1(n7171), .A2(prog_data[5]), .B1(\mem[72][5] ), .B2(n7170), 
        .Z(n3506) );
  OA22D0 U4305 ( .A1(n7171), .A2(prog_data[4]), .B1(\mem[72][4] ), .B2(n7170), 
        .Z(n3505) );
  OA22D0 U4306 ( .A1(n7171), .A2(prog_data[3]), .B1(\mem[72][3] ), .B2(n7170), 
        .Z(n3504) );
  OA22D0 U4307 ( .A1(n7171), .A2(prog_data[2]), .B1(\mem[72][2] ), .B2(n7170), 
        .Z(n3503) );
  OA22D0 U4308 ( .A1(n7171), .A2(prog_data[1]), .B1(\mem[72][1] ), .B2(n7170), 
        .Z(n3502) );
  OA22D0 U4309 ( .A1(n7171), .A2(prog_data[0]), .B1(\mem[72][0] ), .B2(n7170), 
        .Z(n3501) );
  NR2D0 U4310 ( .A1(n7555), .A2(n7184), .ZN(n7172) );
  INVD0 U4311 ( .I(n7172), .ZN(n7173) );
  OA22D0 U4312 ( .A1(n7173), .A2(prog_data[15]), .B1(\mem[73][15] ), .B2(n7172), .Z(n3500) );
  OA22D0 U4313 ( .A1(n7173), .A2(prog_data[14]), .B1(\mem[73][14] ), .B2(n7172), .Z(n3499) );
  OA22D0 U4314 ( .A1(n7173), .A2(prog_data[13]), .B1(\mem[73][13] ), .B2(n7172), .Z(n3498) );
  OA22D0 U4315 ( .A1(n7173), .A2(prog_data[12]), .B1(\mem[73][12] ), .B2(n7172), .Z(n3497) );
  OA22D0 U4316 ( .A1(n7173), .A2(prog_data[11]), .B1(\mem[73][11] ), .B2(n7172), .Z(n3496) );
  OA22D0 U4317 ( .A1(n7173), .A2(prog_data[10]), .B1(\mem[73][10] ), .B2(n7172), .Z(n3495) );
  OA22D0 U4318 ( .A1(n7173), .A2(prog_data[9]), .B1(\mem[73][9] ), .B2(n7172), 
        .Z(n3494) );
  OA22D0 U4319 ( .A1(n7173), .A2(prog_data[8]), .B1(\mem[73][8] ), .B2(n7172), 
        .Z(n3493) );
  OA22D0 U4320 ( .A1(n7173), .A2(prog_data[7]), .B1(\mem[73][7] ), .B2(n7172), 
        .Z(n3492) );
  OA22D0 U4321 ( .A1(n7173), .A2(prog_data[6]), .B1(\mem[73][6] ), .B2(n7172), 
        .Z(n3491) );
  OA22D0 U4322 ( .A1(n7173), .A2(prog_data[5]), .B1(\mem[73][5] ), .B2(n7172), 
        .Z(n3490) );
  OA22D0 U4323 ( .A1(n7173), .A2(prog_data[4]), .B1(\mem[73][4] ), .B2(n7172), 
        .Z(n3489) );
  OA22D0 U4324 ( .A1(n7173), .A2(prog_data[3]), .B1(\mem[73][3] ), .B2(n7172), 
        .Z(n3488) );
  OA22D0 U4325 ( .A1(n7173), .A2(prog_data[2]), .B1(\mem[73][2] ), .B2(n7172), 
        .Z(n3487) );
  OA22D0 U4326 ( .A1(n7173), .A2(prog_data[1]), .B1(\mem[73][1] ), .B2(n7172), 
        .Z(n3486) );
  OA22D0 U4327 ( .A1(n7173), .A2(prog_data[0]), .B1(\mem[73][0] ), .B2(n7172), 
        .Z(n3485) );
  NR2D0 U4328 ( .A1(n7558), .A2(n7184), .ZN(n7174) );
  INVD0 U4329 ( .I(n7174), .ZN(n7175) );
  OA22D0 U4330 ( .A1(n7175), .A2(prog_data[15]), .B1(\mem[74][15] ), .B2(n7174), .Z(n3484) );
  OA22D0 U4331 ( .A1(n7175), .A2(prog_data[14]), .B1(\mem[74][14] ), .B2(n7174), .Z(n3483) );
  OA22D0 U4332 ( .A1(n7175), .A2(prog_data[13]), .B1(\mem[74][13] ), .B2(n7174), .Z(n3482) );
  OA22D0 U4333 ( .A1(n7175), .A2(prog_data[12]), .B1(\mem[74][12] ), .B2(n7174), .Z(n3481) );
  OA22D0 U4334 ( .A1(n7175), .A2(prog_data[11]), .B1(\mem[74][11] ), .B2(n7174), .Z(n3480) );
  OA22D0 U4335 ( .A1(n7175), .A2(prog_data[10]), .B1(\mem[74][10] ), .B2(n7174), .Z(n3479) );
  OA22D0 U4336 ( .A1(n7175), .A2(prog_data[9]), .B1(\mem[74][9] ), .B2(n7174), 
        .Z(n3478) );
  OA22D0 U4337 ( .A1(n7175), .A2(prog_data[8]), .B1(\mem[74][8] ), .B2(n7174), 
        .Z(n3477) );
  OA22D0 U4338 ( .A1(n7175), .A2(prog_data[7]), .B1(\mem[74][7] ), .B2(n7174), 
        .Z(n3476) );
  OA22D0 U4339 ( .A1(n7175), .A2(prog_data[6]), .B1(\mem[74][6] ), .B2(n7174), 
        .Z(n3475) );
  OA22D0 U4340 ( .A1(n7175), .A2(prog_data[5]), .B1(\mem[74][5] ), .B2(n7174), 
        .Z(n3474) );
  OA22D0 U4341 ( .A1(n7175), .A2(prog_data[4]), .B1(\mem[74][4] ), .B2(n7174), 
        .Z(n3473) );
  OA22D0 U4342 ( .A1(n7175), .A2(prog_data[3]), .B1(\mem[74][3] ), .B2(n7174), 
        .Z(n3472) );
  OA22D0 U4343 ( .A1(n7175), .A2(prog_data[2]), .B1(\mem[74][2] ), .B2(n7174), 
        .Z(n3471) );
  OA22D0 U4344 ( .A1(n7175), .A2(prog_data[1]), .B1(\mem[74][1] ), .B2(n7174), 
        .Z(n3470) );
  OA22D0 U4345 ( .A1(n7175), .A2(prog_data[0]), .B1(\mem[74][0] ), .B2(n7174), 
        .Z(n3469) );
  NR2D0 U4346 ( .A1(n7561), .A2(n7184), .ZN(n7176) );
  INVD0 U4347 ( .I(n7176), .ZN(n7177) );
  OA22D0 U4348 ( .A1(n7177), .A2(prog_data[15]), .B1(\mem[75][15] ), .B2(n7176), .Z(n3468) );
  OA22D0 U4349 ( .A1(n7177), .A2(prog_data[14]), .B1(\mem[75][14] ), .B2(n7176), .Z(n3467) );
  OA22D0 U4350 ( .A1(n7177), .A2(prog_data[13]), .B1(\mem[75][13] ), .B2(n7176), .Z(n3466) );
  OA22D0 U4351 ( .A1(n7177), .A2(prog_data[12]), .B1(\mem[75][12] ), .B2(n7176), .Z(n3465) );
  OA22D0 U4352 ( .A1(n7177), .A2(prog_data[11]), .B1(\mem[75][11] ), .B2(n7176), .Z(n3464) );
  OA22D0 U4353 ( .A1(n7177), .A2(prog_data[10]), .B1(\mem[75][10] ), .B2(n7176), .Z(n3463) );
  OA22D0 U4354 ( .A1(n7177), .A2(prog_data[9]), .B1(\mem[75][9] ), .B2(n7176), 
        .Z(n3462) );
  OA22D0 U4355 ( .A1(n7177), .A2(prog_data[8]), .B1(\mem[75][8] ), .B2(n7176), 
        .Z(n3461) );
  OA22D0 U4356 ( .A1(n7177), .A2(prog_data[7]), .B1(\mem[75][7] ), .B2(n7176), 
        .Z(n3460) );
  OA22D0 U4357 ( .A1(n7177), .A2(prog_data[6]), .B1(\mem[75][6] ), .B2(n7176), 
        .Z(n3459) );
  OA22D0 U4358 ( .A1(n7177), .A2(prog_data[5]), .B1(\mem[75][5] ), .B2(n7176), 
        .Z(n3458) );
  OA22D0 U4359 ( .A1(n7177), .A2(prog_data[4]), .B1(\mem[75][4] ), .B2(n7176), 
        .Z(n3457) );
  OA22D0 U4360 ( .A1(n7177), .A2(prog_data[3]), .B1(\mem[75][3] ), .B2(n7176), 
        .Z(n3456) );
  OA22D0 U4361 ( .A1(n7177), .A2(prog_data[2]), .B1(\mem[75][2] ), .B2(n7176), 
        .Z(n3455) );
  OA22D0 U4362 ( .A1(n7177), .A2(prog_data[1]), .B1(\mem[75][1] ), .B2(n7176), 
        .Z(n3454) );
  OA22D0 U4363 ( .A1(n7177), .A2(prog_data[0]), .B1(\mem[75][0] ), .B2(n7176), 
        .Z(n3453) );
  INVD0 U4364 ( .I(n7178), .ZN(n7179) );
  OA22D0 U4365 ( .A1(n7179), .A2(prog_data[15]), .B1(\mem[76][15] ), .B2(n7178), .Z(n3452) );
  OA22D0 U4366 ( .A1(n7179), .A2(prog_data[14]), .B1(\mem[76][14] ), .B2(n7178), .Z(n3451) );
  OA22D0 U4367 ( .A1(n7179), .A2(prog_data[13]), .B1(\mem[76][13] ), .B2(n7178), .Z(n3450) );
  OA22D0 U4368 ( .A1(n7179), .A2(prog_data[12]), .B1(\mem[76][12] ), .B2(n7178), .Z(n3449) );
  OA22D0 U4369 ( .A1(n7179), .A2(prog_data[11]), .B1(\mem[76][11] ), .B2(n7178), .Z(n3448) );
  OA22D0 U4370 ( .A1(n7179), .A2(prog_data[10]), .B1(\mem[76][10] ), .B2(n7178), .Z(n3447) );
  OA22D0 U4371 ( .A1(n7179), .A2(prog_data[9]), .B1(\mem[76][9] ), .B2(n7178), 
        .Z(n3446) );
  OA22D0 U4372 ( .A1(n7179), .A2(prog_data[8]), .B1(\mem[76][8] ), .B2(n7178), 
        .Z(n3445) );
  OA22D0 U4373 ( .A1(n7179), .A2(prog_data[7]), .B1(\mem[76][7] ), .B2(n7178), 
        .Z(n3444) );
  OA22D0 U4374 ( .A1(n7179), .A2(prog_data[6]), .B1(\mem[76][6] ), .B2(n7178), 
        .Z(n3443) );
  OA22D0 U4375 ( .A1(n7179), .A2(prog_data[5]), .B1(\mem[76][5] ), .B2(n7178), 
        .Z(n3442) );
  OA22D0 U4376 ( .A1(n7179), .A2(prog_data[4]), .B1(\mem[76][4] ), .B2(n7178), 
        .Z(n3441) );
  OA22D0 U4377 ( .A1(n7179), .A2(prog_data[3]), .B1(\mem[76][3] ), .B2(n7178), 
        .Z(n3440) );
  OA22D0 U4378 ( .A1(n7179), .A2(prog_data[2]), .B1(\mem[76][2] ), .B2(n7178), 
        .Z(n3439) );
  OA22D0 U4379 ( .A1(n7179), .A2(prog_data[1]), .B1(\mem[76][1] ), .B2(n7178), 
        .Z(n3438) );
  OA22D0 U4380 ( .A1(n7179), .A2(prog_data[0]), .B1(\mem[76][0] ), .B2(n7178), 
        .Z(n3437) );
  NR2D0 U4381 ( .A1(n7567), .A2(n7184), .ZN(n7180) );
  INVD0 U4382 ( .I(n7180), .ZN(n7181) );
  OA22D0 U4383 ( .A1(n7181), .A2(prog_data[15]), .B1(\mem[77][15] ), .B2(n7180), .Z(n3436) );
  OA22D0 U4384 ( .A1(n7181), .A2(prog_data[14]), .B1(\mem[77][14] ), .B2(n7180), .Z(n3435) );
  OA22D0 U4385 ( .A1(n7181), .A2(prog_data[13]), .B1(\mem[77][13] ), .B2(n7180), .Z(n3434) );
  OA22D0 U4386 ( .A1(n7181), .A2(prog_data[12]), .B1(\mem[77][12] ), .B2(n7180), .Z(n3433) );
  OA22D0 U4387 ( .A1(n7181), .A2(prog_data[11]), .B1(\mem[77][11] ), .B2(n7180), .Z(n3432) );
  OA22D0 U4388 ( .A1(n7181), .A2(prog_data[10]), .B1(\mem[77][10] ), .B2(n7180), .Z(n3431) );
  OA22D0 U4389 ( .A1(n7181), .A2(prog_data[9]), .B1(\mem[77][9] ), .B2(n7180), 
        .Z(n3430) );
  OA22D0 U4390 ( .A1(n7181), .A2(prog_data[8]), .B1(\mem[77][8] ), .B2(n7180), 
        .Z(n3429) );
  OA22D0 U4391 ( .A1(n7181), .A2(prog_data[7]), .B1(\mem[77][7] ), .B2(n7180), 
        .Z(n3428) );
  OA22D0 U4392 ( .A1(n7181), .A2(prog_data[6]), .B1(\mem[77][6] ), .B2(n7180), 
        .Z(n3427) );
  OA22D0 U4393 ( .A1(n7181), .A2(prog_data[5]), .B1(\mem[77][5] ), .B2(n7180), 
        .Z(n3426) );
  OA22D0 U4394 ( .A1(n7181), .A2(prog_data[4]), .B1(\mem[77][4] ), .B2(n7180), 
        .Z(n3425) );
  OA22D0 U4395 ( .A1(n7181), .A2(prog_data[3]), .B1(\mem[77][3] ), .B2(n7180), 
        .Z(n3424) );
  OA22D0 U4396 ( .A1(n7181), .A2(prog_data[2]), .B1(\mem[77][2] ), .B2(n7180), 
        .Z(n3423) );
  OA22D0 U4397 ( .A1(n7181), .A2(prog_data[1]), .B1(\mem[77][1] ), .B2(n7180), 
        .Z(n3422) );
  OA22D0 U4398 ( .A1(n7181), .A2(prog_data[0]), .B1(\mem[77][0] ), .B2(n7180), 
        .Z(n3421) );
  NR2D0 U4399 ( .A1(n7570), .A2(n7184), .ZN(n7182) );
  INVD0 U4400 ( .I(n7182), .ZN(n7183) );
  OA22D0 U4401 ( .A1(n7183), .A2(prog_data[15]), .B1(\mem[78][15] ), .B2(n7182), .Z(n3420) );
  OA22D0 U4402 ( .A1(n7183), .A2(prog_data[14]), .B1(\mem[78][14] ), .B2(n7182), .Z(n3419) );
  OA22D0 U4403 ( .A1(n7183), .A2(prog_data[13]), .B1(\mem[78][13] ), .B2(n7182), .Z(n3418) );
  OA22D0 U4404 ( .A1(n7183), .A2(prog_data[12]), .B1(\mem[78][12] ), .B2(n7182), .Z(n3417) );
  OA22D0 U4405 ( .A1(n7183), .A2(prog_data[11]), .B1(\mem[78][11] ), .B2(n7182), .Z(n3416) );
  OA22D0 U4406 ( .A1(n7183), .A2(prog_data[10]), .B1(\mem[78][10] ), .B2(n7182), .Z(n3415) );
  OA22D0 U4407 ( .A1(n7183), .A2(prog_data[9]), .B1(\mem[78][9] ), .B2(n7182), 
        .Z(n3414) );
  OA22D0 U4408 ( .A1(n7183), .A2(prog_data[8]), .B1(\mem[78][8] ), .B2(n7182), 
        .Z(n3413) );
  OA22D0 U4409 ( .A1(n7183), .A2(prog_data[7]), .B1(\mem[78][7] ), .B2(n7182), 
        .Z(n3412) );
  OA22D0 U4410 ( .A1(n7183), .A2(prog_data[6]), .B1(\mem[78][6] ), .B2(n7182), 
        .Z(n3411) );
  OA22D0 U4411 ( .A1(n7183), .A2(prog_data[5]), .B1(\mem[78][5] ), .B2(n7182), 
        .Z(n3410) );
  OA22D0 U4412 ( .A1(n7183), .A2(prog_data[4]), .B1(\mem[78][4] ), .B2(n7182), 
        .Z(n3409) );
  OA22D0 U4413 ( .A1(n7183), .A2(prog_data[3]), .B1(\mem[78][3] ), .B2(n7182), 
        .Z(n3408) );
  OA22D0 U4414 ( .A1(n7183), .A2(prog_data[2]), .B1(\mem[78][2] ), .B2(n7182), 
        .Z(n3407) );
  OA22D0 U4415 ( .A1(n7183), .A2(prog_data[1]), .B1(\mem[78][1] ), .B2(n7182), 
        .Z(n3406) );
  OA22D0 U4416 ( .A1(n7183), .A2(prog_data[0]), .B1(\mem[78][0] ), .B2(n7182), 
        .Z(n3405) );
  NR2D0 U4417 ( .A1(n7574), .A2(n7184), .ZN(n7185) );
  INVD0 U4418 ( .I(n7185), .ZN(n7186) );
  OA22D0 U4419 ( .A1(n7186), .A2(prog_data[15]), .B1(\mem[79][15] ), .B2(n7185), .Z(n3404) );
  OA22D0 U4420 ( .A1(n7186), .A2(prog_data[14]), .B1(\mem[79][14] ), .B2(n7185), .Z(n3403) );
  OA22D0 U4421 ( .A1(n7186), .A2(prog_data[13]), .B1(\mem[79][13] ), .B2(n7185), .Z(n3402) );
  OA22D0 U4422 ( .A1(n7186), .A2(prog_data[12]), .B1(\mem[79][12] ), .B2(n7185), .Z(n3401) );
  OA22D0 U4423 ( .A1(n7186), .A2(prog_data[11]), .B1(\mem[79][11] ), .B2(n7185), .Z(n3400) );
  OA22D0 U4424 ( .A1(n7186), .A2(prog_data[10]), .B1(\mem[79][10] ), .B2(n7185), .Z(n3399) );
  OA22D0 U4425 ( .A1(n7186), .A2(prog_data[9]), .B1(\mem[79][9] ), .B2(n7185), 
        .Z(n3398) );
  OA22D0 U4426 ( .A1(n7186), .A2(prog_data[8]), .B1(\mem[79][8] ), .B2(n7185), 
        .Z(n3397) );
  OA22D0 U4427 ( .A1(n7186), .A2(prog_data[7]), .B1(\mem[79][7] ), .B2(n7185), 
        .Z(n3396) );
  OA22D0 U4428 ( .A1(n7186), .A2(prog_data[6]), .B1(\mem[79][6] ), .B2(n7185), 
        .Z(n3395) );
  OA22D0 U4429 ( .A1(n7186), .A2(prog_data[5]), .B1(\mem[79][5] ), .B2(n7185), 
        .Z(n3394) );
  OA22D0 U4430 ( .A1(n7186), .A2(prog_data[4]), .B1(\mem[79][4] ), .B2(n7185), 
        .Z(n3393) );
  OA22D0 U4431 ( .A1(n7186), .A2(prog_data[3]), .B1(\mem[79][3] ), .B2(n7185), 
        .Z(n3392) );
  OA22D0 U4432 ( .A1(n7186), .A2(prog_data[2]), .B1(\mem[79][2] ), .B2(n7185), 
        .Z(n3391) );
  OA22D0 U4433 ( .A1(n7186), .A2(prog_data[1]), .B1(\mem[79][1] ), .B2(n7185), 
        .Z(n3390) );
  OA22D0 U4434 ( .A1(n7186), .A2(prog_data[0]), .B1(\mem[79][0] ), .B2(n7185), 
        .Z(n3389) );
  ND3D0 U4435 ( .A1(prog_addr[6]), .A2(n7255), .A3(n7187), .ZN(n7218) );
  NR2D0 U4436 ( .A1(n7528), .A2(n7218), .ZN(n7188) );
  INVD0 U4437 ( .I(n7188), .ZN(n7189) );
  OA22D0 U4438 ( .A1(n7189), .A2(prog_data[15]), .B1(\mem[80][15] ), .B2(n7188), .Z(n3388) );
  OA22D0 U4439 ( .A1(n7189), .A2(prog_data[14]), .B1(\mem[80][14] ), .B2(n7188), .Z(n3387) );
  OA22D0 U4440 ( .A1(n7189), .A2(prog_data[13]), .B1(\mem[80][13] ), .B2(n7188), .Z(n3386) );
  OA22D0 U4441 ( .A1(n7189), .A2(prog_data[12]), .B1(\mem[80][12] ), .B2(n7188), .Z(n3385) );
  OA22D0 U4442 ( .A1(n7189), .A2(prog_data[11]), .B1(\mem[80][11] ), .B2(n7188), .Z(n3384) );
  OA22D0 U4443 ( .A1(n7189), .A2(prog_data[10]), .B1(\mem[80][10] ), .B2(n7188), .Z(n3383) );
  OA22D0 U4444 ( .A1(n7189), .A2(prog_data[9]), .B1(\mem[80][9] ), .B2(n7188), 
        .Z(n3382) );
  OA22D0 U4445 ( .A1(n7189), .A2(prog_data[8]), .B1(\mem[80][8] ), .B2(n7188), 
        .Z(n3381) );
  OA22D0 U4446 ( .A1(n7189), .A2(prog_data[7]), .B1(\mem[80][7] ), .B2(n7188), 
        .Z(n3380) );
  OA22D0 U4447 ( .A1(n7189), .A2(prog_data[6]), .B1(\mem[80][6] ), .B2(n7188), 
        .Z(n3379) );
  OA22D0 U4448 ( .A1(n7189), .A2(prog_data[5]), .B1(\mem[80][5] ), .B2(n7188), 
        .Z(n3378) );
  OA22D0 U4449 ( .A1(n7189), .A2(prog_data[4]), .B1(\mem[80][4] ), .B2(n7188), 
        .Z(n3377) );
  OA22D0 U4450 ( .A1(n7189), .A2(prog_data[3]), .B1(\mem[80][3] ), .B2(n7188), 
        .Z(n3376) );
  OA22D0 U4451 ( .A1(n7189), .A2(prog_data[2]), .B1(\mem[80][2] ), .B2(n7188), 
        .Z(n3375) );
  OA22D0 U4452 ( .A1(n7189), .A2(prog_data[1]), .B1(\mem[80][1] ), .B2(n7188), 
        .Z(n3374) );
  OA22D0 U4453 ( .A1(n7189), .A2(prog_data[0]), .B1(\mem[80][0] ), .B2(n7188), 
        .Z(n3373) );
  NR2D0 U4454 ( .A1(n7531), .A2(n7218), .ZN(n7190) );
  INVD0 U4455 ( .I(n7190), .ZN(n7191) );
  OA22D0 U4456 ( .A1(n7191), .A2(prog_data[15]), .B1(\mem[81][15] ), .B2(n7190), .Z(n3372) );
  OA22D0 U4457 ( .A1(n7191), .A2(prog_data[14]), .B1(\mem[81][14] ), .B2(n7190), .Z(n3371) );
  OA22D0 U4458 ( .A1(n7191), .A2(prog_data[13]), .B1(\mem[81][13] ), .B2(n7190), .Z(n3370) );
  OA22D0 U4459 ( .A1(n7191), .A2(prog_data[12]), .B1(\mem[81][12] ), .B2(n7190), .Z(n3369) );
  OA22D0 U4460 ( .A1(n7191), .A2(prog_data[11]), .B1(\mem[81][11] ), .B2(n7190), .Z(n3368) );
  OA22D0 U4461 ( .A1(n7191), .A2(prog_data[10]), .B1(\mem[81][10] ), .B2(n7190), .Z(n3367) );
  OA22D0 U4462 ( .A1(n7191), .A2(prog_data[9]), .B1(\mem[81][9] ), .B2(n7190), 
        .Z(n3366) );
  OA22D0 U4463 ( .A1(n7191), .A2(prog_data[8]), .B1(\mem[81][8] ), .B2(n7190), 
        .Z(n3365) );
  OA22D0 U4464 ( .A1(n7191), .A2(prog_data[7]), .B1(\mem[81][7] ), .B2(n7190), 
        .Z(n3364) );
  OA22D0 U4465 ( .A1(n7191), .A2(prog_data[6]), .B1(\mem[81][6] ), .B2(n7190), 
        .Z(n3363) );
  OA22D0 U4466 ( .A1(n7191), .A2(prog_data[5]), .B1(\mem[81][5] ), .B2(n7190), 
        .Z(n3362) );
  OA22D0 U4467 ( .A1(n7191), .A2(prog_data[4]), .B1(\mem[81][4] ), .B2(n7190), 
        .Z(n3361) );
  OA22D0 U4468 ( .A1(n7191), .A2(prog_data[3]), .B1(\mem[81][3] ), .B2(n7190), 
        .Z(n3360) );
  OA22D0 U4469 ( .A1(n7191), .A2(prog_data[2]), .B1(\mem[81][2] ), .B2(n7190), 
        .Z(n3359) );
  OA22D0 U4470 ( .A1(n7191), .A2(prog_data[1]), .B1(\mem[81][1] ), .B2(n7190), 
        .Z(n3358) );
  OA22D0 U4471 ( .A1(n7191), .A2(prog_data[0]), .B1(\mem[81][0] ), .B2(n7190), 
        .Z(n3357) );
  NR2D0 U4472 ( .A1(n7534), .A2(n7218), .ZN(n7192) );
  INVD0 U4473 ( .I(n7192), .ZN(n7193) );
  OA22D0 U4474 ( .A1(n7193), .A2(prog_data[15]), .B1(\mem[82][15] ), .B2(n7192), .Z(n3356) );
  OA22D0 U4475 ( .A1(n7193), .A2(prog_data[14]), .B1(\mem[82][14] ), .B2(n7192), .Z(n3355) );
  OA22D0 U4476 ( .A1(n7193), .A2(prog_data[13]), .B1(\mem[82][13] ), .B2(n7192), .Z(n3354) );
  OA22D0 U4477 ( .A1(n7193), .A2(prog_data[12]), .B1(\mem[82][12] ), .B2(n7192), .Z(n3353) );
  OA22D0 U4478 ( .A1(n7193), .A2(prog_data[11]), .B1(\mem[82][11] ), .B2(n7192), .Z(n3352) );
  OA22D0 U4479 ( .A1(n7193), .A2(prog_data[10]), .B1(\mem[82][10] ), .B2(n7192), .Z(n3351) );
  OA22D0 U4480 ( .A1(n7193), .A2(prog_data[9]), .B1(\mem[82][9] ), .B2(n7192), 
        .Z(n3350) );
  OA22D0 U4481 ( .A1(n7193), .A2(prog_data[8]), .B1(\mem[82][8] ), .B2(n7192), 
        .Z(n3349) );
  OA22D0 U4482 ( .A1(n7193), .A2(prog_data[7]), .B1(\mem[82][7] ), .B2(n7192), 
        .Z(n3348) );
  OA22D0 U4483 ( .A1(n7193), .A2(prog_data[6]), .B1(\mem[82][6] ), .B2(n7192), 
        .Z(n3347) );
  OA22D0 U4484 ( .A1(n7193), .A2(prog_data[5]), .B1(\mem[82][5] ), .B2(n7192), 
        .Z(n3346) );
  OA22D0 U4485 ( .A1(n7193), .A2(prog_data[4]), .B1(\mem[82][4] ), .B2(n7192), 
        .Z(n3345) );
  OA22D0 U4486 ( .A1(n7193), .A2(prog_data[3]), .B1(\mem[82][3] ), .B2(n7192), 
        .Z(n3344) );
  OA22D0 U4487 ( .A1(n7193), .A2(prog_data[2]), .B1(\mem[82][2] ), .B2(n7192), 
        .Z(n3343) );
  OA22D0 U4488 ( .A1(n7193), .A2(prog_data[1]), .B1(\mem[82][1] ), .B2(n7192), 
        .Z(n3342) );
  OA22D0 U4489 ( .A1(n7193), .A2(prog_data[0]), .B1(\mem[82][0] ), .B2(n7192), 
        .Z(n3341) );
  NR2D0 U4490 ( .A1(n7537), .A2(n7218), .ZN(n7194) );
  INVD0 U4491 ( .I(n7194), .ZN(n7195) );
  OA22D0 U4492 ( .A1(n7195), .A2(prog_data[15]), .B1(\mem[83][15] ), .B2(n7194), .Z(n3340) );
  OA22D0 U4493 ( .A1(n7195), .A2(prog_data[14]), .B1(\mem[83][14] ), .B2(n7194), .Z(n3339) );
  OA22D0 U4494 ( .A1(n7195), .A2(prog_data[13]), .B1(\mem[83][13] ), .B2(n7194), .Z(n3338) );
  OA22D0 U4495 ( .A1(n7195), .A2(prog_data[12]), .B1(\mem[83][12] ), .B2(n7194), .Z(n3337) );
  OA22D0 U4496 ( .A1(n7195), .A2(prog_data[11]), .B1(\mem[83][11] ), .B2(n7194), .Z(n3336) );
  OA22D0 U4497 ( .A1(n7195), .A2(prog_data[10]), .B1(\mem[83][10] ), .B2(n7194), .Z(n3335) );
  OA22D0 U4498 ( .A1(n7195), .A2(prog_data[9]), .B1(\mem[83][9] ), .B2(n7194), 
        .Z(n3334) );
  OA22D0 U4499 ( .A1(n7195), .A2(prog_data[8]), .B1(\mem[83][8] ), .B2(n7194), 
        .Z(n3333) );
  OA22D0 U4500 ( .A1(n7195), .A2(prog_data[7]), .B1(\mem[83][7] ), .B2(n7194), 
        .Z(n3332) );
  OA22D0 U4501 ( .A1(n7195), .A2(prog_data[6]), .B1(\mem[83][6] ), .B2(n7194), 
        .Z(n3331) );
  OA22D0 U4502 ( .A1(n7195), .A2(prog_data[5]), .B1(\mem[83][5] ), .B2(n7194), 
        .Z(n3330) );
  OA22D0 U4503 ( .A1(n7195), .A2(prog_data[4]), .B1(\mem[83][4] ), .B2(n7194), 
        .Z(n3329) );
  OA22D0 U4504 ( .A1(n7195), .A2(prog_data[3]), .B1(\mem[83][3] ), .B2(n7194), 
        .Z(n3328) );
  OA22D0 U4505 ( .A1(n7195), .A2(prog_data[2]), .B1(\mem[83][2] ), .B2(n7194), 
        .Z(n3327) );
  OA22D0 U4506 ( .A1(n7195), .A2(prog_data[1]), .B1(\mem[83][1] ), .B2(n7194), 
        .Z(n3326) );
  OA22D0 U4507 ( .A1(n7195), .A2(prog_data[0]), .B1(\mem[83][0] ), .B2(n7194), 
        .Z(n3325) );
  NR2D0 U4508 ( .A1(n7540), .A2(n7218), .ZN(n7196) );
  OA22D0 U4509 ( .A1(n7197), .A2(prog_data[15]), .B1(\mem[84][15] ), .B2(n7196), .Z(n3324) );
  OA22D0 U4510 ( .A1(n7197), .A2(prog_data[14]), .B1(\mem[84][14] ), .B2(n7196), .Z(n3323) );
  OA22D0 U4511 ( .A1(n7197), .A2(prog_data[13]), .B1(\mem[84][13] ), .B2(n7196), .Z(n3322) );
  OA22D0 U4512 ( .A1(n7197), .A2(prog_data[12]), .B1(\mem[84][12] ), .B2(n7196), .Z(n3321) );
  OA22D0 U4513 ( .A1(n7197), .A2(prog_data[11]), .B1(\mem[84][11] ), .B2(n7196), .Z(n3320) );
  OA22D0 U4514 ( .A1(n7197), .A2(prog_data[10]), .B1(\mem[84][10] ), .B2(n7196), .Z(n3319) );
  OA22D0 U4515 ( .A1(n7197), .A2(prog_data[9]), .B1(\mem[84][9] ), .B2(n7196), 
        .Z(n3318) );
  OA22D0 U4516 ( .A1(n7197), .A2(prog_data[8]), .B1(\mem[84][8] ), .B2(n7196), 
        .Z(n3317) );
  OA22D0 U4517 ( .A1(n7197), .A2(prog_data[7]), .B1(\mem[84][7] ), .B2(n7196), 
        .Z(n3316) );
  OA22D0 U4518 ( .A1(n7197), .A2(prog_data[6]), .B1(\mem[84][6] ), .B2(n7196), 
        .Z(n3315) );
  OA22D0 U4519 ( .A1(n7197), .A2(prog_data[5]), .B1(\mem[84][5] ), .B2(n7196), 
        .Z(n3314) );
  OA22D0 U4520 ( .A1(n7197), .A2(prog_data[4]), .B1(\mem[84][4] ), .B2(n7196), 
        .Z(n3313) );
  OA22D0 U4521 ( .A1(n7197), .A2(prog_data[3]), .B1(\mem[84][3] ), .B2(n7196), 
        .Z(n3312) );
  OA22D0 U4522 ( .A1(n7197), .A2(prog_data[2]), .B1(\mem[84][2] ), .B2(n7196), 
        .Z(n3311) );
  OA22D0 U4523 ( .A1(n7197), .A2(prog_data[1]), .B1(\mem[84][1] ), .B2(n7196), 
        .Z(n3310) );
  OA22D0 U4524 ( .A1(n7197), .A2(prog_data[0]), .B1(\mem[84][0] ), .B2(n7196), 
        .Z(n3309) );
  NR2D0 U4525 ( .A1(n7543), .A2(n7218), .ZN(n7198) );
  INVD0 U4526 ( .I(n7198), .ZN(n7199) );
  OA22D0 U4527 ( .A1(n7199), .A2(prog_data[15]), .B1(\mem[85][15] ), .B2(n7198), .Z(n3308) );
  OA22D0 U4528 ( .A1(n7199), .A2(prog_data[14]), .B1(\mem[85][14] ), .B2(n7198), .Z(n3307) );
  OA22D0 U4529 ( .A1(n7199), .A2(prog_data[13]), .B1(\mem[85][13] ), .B2(n7198), .Z(n3306) );
  OA22D0 U4530 ( .A1(n7199), .A2(prog_data[12]), .B1(\mem[85][12] ), .B2(n7198), .Z(n3305) );
  OA22D0 U4531 ( .A1(n7199), .A2(prog_data[11]), .B1(\mem[85][11] ), .B2(n7198), .Z(n3304) );
  OA22D0 U4532 ( .A1(n7199), .A2(prog_data[10]), .B1(\mem[85][10] ), .B2(n7198), .Z(n3303) );
  OA22D0 U4533 ( .A1(n7199), .A2(prog_data[9]), .B1(\mem[85][9] ), .B2(n7198), 
        .Z(n3302) );
  OA22D0 U4534 ( .A1(n7199), .A2(prog_data[8]), .B1(\mem[85][8] ), .B2(n7198), 
        .Z(n3301) );
  OA22D0 U4535 ( .A1(n7199), .A2(prog_data[7]), .B1(\mem[85][7] ), .B2(n7198), 
        .Z(n3300) );
  OA22D0 U4536 ( .A1(n7199), .A2(prog_data[6]), .B1(\mem[85][6] ), .B2(n7198), 
        .Z(n3299) );
  OA22D0 U4537 ( .A1(n7199), .A2(prog_data[5]), .B1(\mem[85][5] ), .B2(n7198), 
        .Z(n3298) );
  OA22D0 U4538 ( .A1(n7199), .A2(prog_data[4]), .B1(\mem[85][4] ), .B2(n7198), 
        .Z(n3297) );
  OA22D0 U4539 ( .A1(n7199), .A2(prog_data[3]), .B1(\mem[85][3] ), .B2(n7198), 
        .Z(n3296) );
  OA22D0 U4540 ( .A1(n7199), .A2(prog_data[2]), .B1(\mem[85][2] ), .B2(n7198), 
        .Z(n3295) );
  OA22D0 U4541 ( .A1(n7199), .A2(prog_data[1]), .B1(\mem[85][1] ), .B2(n7198), 
        .Z(n3294) );
  OA22D0 U4542 ( .A1(n7199), .A2(prog_data[0]), .B1(\mem[85][0] ), .B2(n7198), 
        .Z(n3293) );
  NR2D0 U4543 ( .A1(n7546), .A2(n7218), .ZN(n7200) );
  INVD0 U4544 ( .I(n7200), .ZN(n7201) );
  OA22D0 U4545 ( .A1(n7201), .A2(prog_data[15]), .B1(\mem[86][15] ), .B2(n7200), .Z(n3292) );
  OA22D0 U4546 ( .A1(n7201), .A2(prog_data[14]), .B1(\mem[86][14] ), .B2(n7200), .Z(n3291) );
  OA22D0 U4547 ( .A1(n7201), .A2(prog_data[13]), .B1(\mem[86][13] ), .B2(n7200), .Z(n3290) );
  OA22D0 U4548 ( .A1(n7201), .A2(prog_data[12]), .B1(\mem[86][12] ), .B2(n7200), .Z(n3289) );
  OA22D0 U4549 ( .A1(n7201), .A2(prog_data[11]), .B1(\mem[86][11] ), .B2(n7200), .Z(n3288) );
  OA22D0 U4550 ( .A1(n7201), .A2(prog_data[10]), .B1(\mem[86][10] ), .B2(n7200), .Z(n3287) );
  OA22D0 U4551 ( .A1(n7201), .A2(prog_data[9]), .B1(\mem[86][9] ), .B2(n7200), 
        .Z(n3286) );
  OA22D0 U4552 ( .A1(n7201), .A2(prog_data[8]), .B1(\mem[86][8] ), .B2(n7200), 
        .Z(n3285) );
  OA22D0 U4553 ( .A1(n7201), .A2(prog_data[7]), .B1(\mem[86][7] ), .B2(n7200), 
        .Z(n3284) );
  OA22D0 U4554 ( .A1(n7201), .A2(prog_data[6]), .B1(\mem[86][6] ), .B2(n7200), 
        .Z(n3283) );
  OA22D0 U4555 ( .A1(n7201), .A2(prog_data[5]), .B1(\mem[86][5] ), .B2(n7200), 
        .Z(n3282) );
  OA22D0 U4556 ( .A1(n7201), .A2(prog_data[4]), .B1(\mem[86][4] ), .B2(n7200), 
        .Z(n3281) );
  OA22D0 U4557 ( .A1(n7201), .A2(prog_data[3]), .B1(\mem[86][3] ), .B2(n7200), 
        .Z(n3280) );
  OA22D0 U4558 ( .A1(n7201), .A2(prog_data[2]), .B1(\mem[86][2] ), .B2(n7200), 
        .Z(n3279) );
  OA22D0 U4559 ( .A1(n7201), .A2(prog_data[1]), .B1(\mem[86][1] ), .B2(n7200), 
        .Z(n3278) );
  OA22D0 U4560 ( .A1(n7201), .A2(prog_data[0]), .B1(\mem[86][0] ), .B2(n7200), 
        .Z(n3277) );
  NR2D0 U4561 ( .A1(n7549), .A2(n7218), .ZN(n7202) );
  INVD0 U4562 ( .I(n7202), .ZN(n7203) );
  OA22D0 U4563 ( .A1(n7203), .A2(prog_data[15]), .B1(\mem[87][15] ), .B2(n7202), .Z(n3276) );
  OA22D0 U4564 ( .A1(n7203), .A2(prog_data[14]), .B1(\mem[87][14] ), .B2(n7202), .Z(n3275) );
  OA22D0 U4565 ( .A1(n7203), .A2(prog_data[13]), .B1(\mem[87][13] ), .B2(n7202), .Z(n3274) );
  OA22D0 U4566 ( .A1(n7203), .A2(prog_data[12]), .B1(\mem[87][12] ), .B2(n7202), .Z(n3273) );
  OA22D0 U4567 ( .A1(n7203), .A2(prog_data[11]), .B1(\mem[87][11] ), .B2(n7202), .Z(n3272) );
  OA22D0 U4568 ( .A1(n7203), .A2(prog_data[10]), .B1(\mem[87][10] ), .B2(n7202), .Z(n3271) );
  OA22D0 U4569 ( .A1(n7203), .A2(prog_data[9]), .B1(\mem[87][9] ), .B2(n7202), 
        .Z(n3270) );
  OA22D0 U4570 ( .A1(n7203), .A2(prog_data[8]), .B1(\mem[87][8] ), .B2(n7202), 
        .Z(n3269) );
  OA22D0 U4571 ( .A1(n7203), .A2(prog_data[7]), .B1(\mem[87][7] ), .B2(n7202), 
        .Z(n3268) );
  OA22D0 U4572 ( .A1(n7203), .A2(prog_data[6]), .B1(\mem[87][6] ), .B2(n7202), 
        .Z(n3267) );
  OA22D0 U4573 ( .A1(n7203), .A2(prog_data[5]), .B1(\mem[87][5] ), .B2(n7202), 
        .Z(n3266) );
  OA22D0 U4574 ( .A1(n7203), .A2(prog_data[4]), .B1(\mem[87][4] ), .B2(n7202), 
        .Z(n3265) );
  OA22D0 U4575 ( .A1(n7203), .A2(prog_data[3]), .B1(\mem[87][3] ), .B2(n7202), 
        .Z(n3264) );
  OA22D0 U4576 ( .A1(n7203), .A2(prog_data[2]), .B1(\mem[87][2] ), .B2(n7202), 
        .Z(n3263) );
  OA22D0 U4577 ( .A1(n7203), .A2(prog_data[1]), .B1(\mem[87][1] ), .B2(n7202), 
        .Z(n3262) );
  OA22D0 U4578 ( .A1(n7203), .A2(prog_data[0]), .B1(\mem[87][0] ), .B2(n7202), 
        .Z(n3261) );
  NR2D0 U4579 ( .A1(n7552), .A2(n7218), .ZN(n7204) );
  INVD0 U4580 ( .I(n7204), .ZN(n7205) );
  OA22D0 U4581 ( .A1(n7205), .A2(prog_data[15]), .B1(\mem[88][15] ), .B2(n7204), .Z(n3260) );
  OA22D0 U4582 ( .A1(n7205), .A2(prog_data[14]), .B1(\mem[88][14] ), .B2(n7204), .Z(n3259) );
  OA22D0 U4583 ( .A1(n7205), .A2(prog_data[13]), .B1(\mem[88][13] ), .B2(n7204), .Z(n3258) );
  OA22D0 U4584 ( .A1(n7205), .A2(prog_data[12]), .B1(\mem[88][12] ), .B2(n7204), .Z(n3257) );
  OA22D0 U4585 ( .A1(n7205), .A2(prog_data[11]), .B1(\mem[88][11] ), .B2(n7204), .Z(n3256) );
  OA22D0 U4586 ( .A1(n7205), .A2(prog_data[10]), .B1(\mem[88][10] ), .B2(n7204), .Z(n3255) );
  OA22D0 U4587 ( .A1(n7205), .A2(prog_data[9]), .B1(\mem[88][9] ), .B2(n7204), 
        .Z(n3254) );
  OA22D0 U4588 ( .A1(n7205), .A2(prog_data[8]), .B1(\mem[88][8] ), .B2(n7204), 
        .Z(n3253) );
  OA22D0 U4589 ( .A1(n7205), .A2(prog_data[7]), .B1(\mem[88][7] ), .B2(n7204), 
        .Z(n3252) );
  OA22D0 U4590 ( .A1(n7205), .A2(prog_data[6]), .B1(\mem[88][6] ), .B2(n7204), 
        .Z(n3251) );
  OA22D0 U4591 ( .A1(n7205), .A2(prog_data[5]), .B1(\mem[88][5] ), .B2(n7204), 
        .Z(n3250) );
  OA22D0 U4592 ( .A1(n7205), .A2(prog_data[4]), .B1(\mem[88][4] ), .B2(n7204), 
        .Z(n3249) );
  OA22D0 U4593 ( .A1(n7205), .A2(prog_data[3]), .B1(\mem[88][3] ), .B2(n7204), 
        .Z(n3248) );
  OA22D0 U4594 ( .A1(n7205), .A2(prog_data[2]), .B1(\mem[88][2] ), .B2(n7204), 
        .Z(n3247) );
  OA22D0 U4595 ( .A1(n7205), .A2(prog_data[1]), .B1(\mem[88][1] ), .B2(n7204), 
        .Z(n3246) );
  OA22D0 U4596 ( .A1(n7205), .A2(prog_data[0]), .B1(\mem[88][0] ), .B2(n7204), 
        .Z(n3245) );
  NR2D0 U4597 ( .A1(n7555), .A2(n7218), .ZN(n7206) );
  INVD0 U4598 ( .I(n7206), .ZN(n7207) );
  OA22D0 U4599 ( .A1(n7207), .A2(prog_data[15]), .B1(\mem[89][15] ), .B2(n7206), .Z(n3244) );
  OA22D0 U4600 ( .A1(n7207), .A2(prog_data[14]), .B1(\mem[89][14] ), .B2(n7206), .Z(n3243) );
  OA22D0 U4601 ( .A1(n7207), .A2(prog_data[13]), .B1(\mem[89][13] ), .B2(n7206), .Z(n3242) );
  OA22D0 U4602 ( .A1(n7207), .A2(prog_data[12]), .B1(\mem[89][12] ), .B2(n7206), .Z(n3241) );
  OA22D0 U4603 ( .A1(n7207), .A2(prog_data[11]), .B1(\mem[89][11] ), .B2(n7206), .Z(n3240) );
  OA22D0 U4604 ( .A1(n7207), .A2(prog_data[10]), .B1(\mem[89][10] ), .B2(n7206), .Z(n3239) );
  OA22D0 U4605 ( .A1(n7207), .A2(prog_data[9]), .B1(\mem[89][9] ), .B2(n7206), 
        .Z(n3238) );
  OA22D0 U4606 ( .A1(n7207), .A2(prog_data[8]), .B1(\mem[89][8] ), .B2(n7206), 
        .Z(n3237) );
  OA22D0 U4607 ( .A1(n7207), .A2(prog_data[7]), .B1(\mem[89][7] ), .B2(n7206), 
        .Z(n3236) );
  OA22D0 U4608 ( .A1(n7207), .A2(prog_data[6]), .B1(\mem[89][6] ), .B2(n7206), 
        .Z(n3235) );
  OA22D0 U4609 ( .A1(n7207), .A2(prog_data[5]), .B1(\mem[89][5] ), .B2(n7206), 
        .Z(n3234) );
  OA22D0 U4610 ( .A1(n7207), .A2(prog_data[4]), .B1(\mem[89][4] ), .B2(n7206), 
        .Z(n3233) );
  OA22D0 U4611 ( .A1(n7207), .A2(prog_data[3]), .B1(\mem[89][3] ), .B2(n7206), 
        .Z(n3232) );
  OA22D0 U4612 ( .A1(n7207), .A2(prog_data[2]), .B1(\mem[89][2] ), .B2(n7206), 
        .Z(n3231) );
  OA22D0 U4613 ( .A1(n7207), .A2(prog_data[1]), .B1(\mem[89][1] ), .B2(n7206), 
        .Z(n3230) );
  OA22D0 U4614 ( .A1(n7207), .A2(prog_data[0]), .B1(\mem[89][0] ), .B2(n7206), 
        .Z(n3229) );
  NR2D0 U4615 ( .A1(n7558), .A2(n7218), .ZN(n7208) );
  INVD0 U4616 ( .I(n7208), .ZN(n7209) );
  OA22D0 U4617 ( .A1(n7209), .A2(prog_data[15]), .B1(\mem[90][15] ), .B2(n7208), .Z(n3228) );
  OA22D0 U4618 ( .A1(n7209), .A2(prog_data[14]), .B1(\mem[90][14] ), .B2(n7208), .Z(n3227) );
  OA22D0 U4619 ( .A1(n7209), .A2(prog_data[13]), .B1(\mem[90][13] ), .B2(n7208), .Z(n3226) );
  OA22D0 U4620 ( .A1(n7209), .A2(prog_data[12]), .B1(\mem[90][12] ), .B2(n7208), .Z(n3225) );
  OA22D0 U4621 ( .A1(n7209), .A2(prog_data[11]), .B1(\mem[90][11] ), .B2(n7208), .Z(n3224) );
  OA22D0 U4622 ( .A1(n7209), .A2(prog_data[10]), .B1(\mem[90][10] ), .B2(n7208), .Z(n3223) );
  OA22D0 U4623 ( .A1(n7209), .A2(prog_data[9]), .B1(\mem[90][9] ), .B2(n7208), 
        .Z(n3222) );
  OA22D0 U4624 ( .A1(n7209), .A2(prog_data[8]), .B1(\mem[90][8] ), .B2(n7208), 
        .Z(n3221) );
  OA22D0 U4625 ( .A1(n7209), .A2(prog_data[7]), .B1(\mem[90][7] ), .B2(n7208), 
        .Z(n3220) );
  OA22D0 U4626 ( .A1(n7209), .A2(prog_data[6]), .B1(\mem[90][6] ), .B2(n7208), 
        .Z(n3219) );
  OA22D0 U4627 ( .A1(n7209), .A2(prog_data[5]), .B1(\mem[90][5] ), .B2(n7208), 
        .Z(n3218) );
  OA22D0 U4628 ( .A1(n7209), .A2(prog_data[4]), .B1(\mem[90][4] ), .B2(n7208), 
        .Z(n3217) );
  OA22D0 U4629 ( .A1(n7209), .A2(prog_data[3]), .B1(\mem[90][3] ), .B2(n7208), 
        .Z(n3216) );
  OA22D0 U4630 ( .A1(n7209), .A2(prog_data[2]), .B1(\mem[90][2] ), .B2(n7208), 
        .Z(n3215) );
  OA22D0 U4631 ( .A1(n7209), .A2(prog_data[1]), .B1(\mem[90][1] ), .B2(n7208), 
        .Z(n3214) );
  OA22D0 U4632 ( .A1(n7209), .A2(prog_data[0]), .B1(\mem[90][0] ), .B2(n7208), 
        .Z(n3213) );
  INVD0 U4633 ( .I(n7210), .ZN(n7211) );
  OA22D0 U4634 ( .A1(n7211), .A2(prog_data[15]), .B1(\mem[91][15] ), .B2(n7210), .Z(n3212) );
  OA22D0 U4635 ( .A1(n7211), .A2(prog_data[14]), .B1(\mem[91][14] ), .B2(n7210), .Z(n3211) );
  OA22D0 U4636 ( .A1(n7211), .A2(prog_data[13]), .B1(\mem[91][13] ), .B2(n7210), .Z(n3210) );
  OA22D0 U4637 ( .A1(n7211), .A2(prog_data[12]), .B1(\mem[91][12] ), .B2(n7210), .Z(n3209) );
  OA22D0 U4638 ( .A1(n7211), .A2(prog_data[11]), .B1(\mem[91][11] ), .B2(n7210), .Z(n3208) );
  OA22D0 U4639 ( .A1(n7211), .A2(prog_data[10]), .B1(\mem[91][10] ), .B2(n7210), .Z(n3207) );
  OA22D0 U4640 ( .A1(n7211), .A2(prog_data[9]), .B1(\mem[91][9] ), .B2(n7210), 
        .Z(n3206) );
  OA22D0 U4641 ( .A1(n7211), .A2(prog_data[8]), .B1(\mem[91][8] ), .B2(n7210), 
        .Z(n3205) );
  OA22D0 U4642 ( .A1(n7211), .A2(prog_data[7]), .B1(\mem[91][7] ), .B2(n7210), 
        .Z(n3204) );
  OA22D0 U4643 ( .A1(n7211), .A2(prog_data[6]), .B1(\mem[91][6] ), .B2(n7210), 
        .Z(n3203) );
  OA22D0 U4644 ( .A1(n7211), .A2(prog_data[5]), .B1(\mem[91][5] ), .B2(n7210), 
        .Z(n3202) );
  OA22D0 U4645 ( .A1(n7211), .A2(prog_data[4]), .B1(\mem[91][4] ), .B2(n7210), 
        .Z(n3201) );
  OA22D0 U4646 ( .A1(n7211), .A2(prog_data[3]), .B1(\mem[91][3] ), .B2(n7210), 
        .Z(n3200) );
  OA22D0 U4647 ( .A1(n7211), .A2(prog_data[2]), .B1(\mem[91][2] ), .B2(n7210), 
        .Z(n3199) );
  OA22D0 U4648 ( .A1(n7211), .A2(prog_data[1]), .B1(\mem[91][1] ), .B2(n7210), 
        .Z(n3198) );
  OA22D0 U4649 ( .A1(n7211), .A2(prog_data[0]), .B1(\mem[91][0] ), .B2(n7210), 
        .Z(n3197) );
  NR2D0 U4650 ( .A1(n7564), .A2(n7218), .ZN(n7212) );
  INVD0 U4651 ( .I(n7212), .ZN(n7213) );
  OA22D0 U4652 ( .A1(n7213), .A2(prog_data[15]), .B1(\mem[92][15] ), .B2(n7212), .Z(n3196) );
  OA22D0 U4653 ( .A1(n7213), .A2(prog_data[14]), .B1(\mem[92][14] ), .B2(n7212), .Z(n3195) );
  OA22D0 U4654 ( .A1(n7213), .A2(prog_data[13]), .B1(\mem[92][13] ), .B2(n7212), .Z(n3194) );
  OA22D0 U4655 ( .A1(n7213), .A2(prog_data[12]), .B1(\mem[92][12] ), .B2(n7212), .Z(n3193) );
  OA22D0 U4656 ( .A1(n7213), .A2(prog_data[11]), .B1(\mem[92][11] ), .B2(n7212), .Z(n3192) );
  OA22D0 U4657 ( .A1(n7213), .A2(prog_data[10]), .B1(\mem[92][10] ), .B2(n7212), .Z(n3191) );
  OA22D0 U4658 ( .A1(n7213), .A2(prog_data[9]), .B1(\mem[92][9] ), .B2(n7212), 
        .Z(n3190) );
  OA22D0 U4659 ( .A1(n7213), .A2(prog_data[8]), .B1(\mem[92][8] ), .B2(n7212), 
        .Z(n3189) );
  OA22D0 U4660 ( .A1(n7213), .A2(prog_data[7]), .B1(\mem[92][7] ), .B2(n7212), 
        .Z(n3188) );
  OA22D0 U4661 ( .A1(n7213), .A2(prog_data[6]), .B1(\mem[92][6] ), .B2(n7212), 
        .Z(n3187) );
  OA22D0 U4662 ( .A1(n7213), .A2(prog_data[5]), .B1(\mem[92][5] ), .B2(n7212), 
        .Z(n3186) );
  OA22D0 U4663 ( .A1(n7213), .A2(prog_data[4]), .B1(\mem[92][4] ), .B2(n7212), 
        .Z(n3185) );
  OA22D0 U4664 ( .A1(n7213), .A2(prog_data[3]), .B1(\mem[92][3] ), .B2(n7212), 
        .Z(n3184) );
  OA22D0 U4665 ( .A1(n7213), .A2(prog_data[2]), .B1(\mem[92][2] ), .B2(n7212), 
        .Z(n3183) );
  OA22D0 U4666 ( .A1(n7213), .A2(prog_data[1]), .B1(\mem[92][1] ), .B2(n7212), 
        .Z(n3182) );
  OA22D0 U4667 ( .A1(n7213), .A2(prog_data[0]), .B1(\mem[92][0] ), .B2(n7212), 
        .Z(n3181) );
  NR2D0 U4668 ( .A1(n7567), .A2(n7218), .ZN(n7214) );
  INVD0 U4669 ( .I(n7214), .ZN(n7215) );
  OA22D0 U4670 ( .A1(n7215), .A2(prog_data[15]), .B1(\mem[93][15] ), .B2(n7214), .Z(n3180) );
  OA22D0 U4671 ( .A1(n7215), .A2(prog_data[14]), .B1(\mem[93][14] ), .B2(n7214), .Z(n3179) );
  OA22D0 U4672 ( .A1(n7215), .A2(prog_data[13]), .B1(\mem[93][13] ), .B2(n7214), .Z(n3178) );
  OA22D0 U4673 ( .A1(n7215), .A2(prog_data[12]), .B1(\mem[93][12] ), .B2(n7214), .Z(n3177) );
  OA22D0 U4674 ( .A1(n7215), .A2(prog_data[11]), .B1(\mem[93][11] ), .B2(n7214), .Z(n3176) );
  OA22D0 U4675 ( .A1(n7215), .A2(prog_data[10]), .B1(\mem[93][10] ), .B2(n7214), .Z(n3175) );
  OA22D0 U4676 ( .A1(n7215), .A2(prog_data[9]), .B1(\mem[93][9] ), .B2(n7214), 
        .Z(n3174) );
  OA22D0 U4677 ( .A1(n7215), .A2(prog_data[8]), .B1(\mem[93][8] ), .B2(n7214), 
        .Z(n3173) );
  OA22D0 U4678 ( .A1(n7215), .A2(prog_data[7]), .B1(\mem[93][7] ), .B2(n7214), 
        .Z(n3172) );
  OA22D0 U4679 ( .A1(n7215), .A2(prog_data[6]), .B1(\mem[93][6] ), .B2(n7214), 
        .Z(n3171) );
  OA22D0 U4680 ( .A1(n7215), .A2(prog_data[5]), .B1(\mem[93][5] ), .B2(n7214), 
        .Z(n3170) );
  OA22D0 U4681 ( .A1(n7215), .A2(prog_data[4]), .B1(\mem[93][4] ), .B2(n7214), 
        .Z(n3169) );
  OA22D0 U4682 ( .A1(n7215), .A2(prog_data[3]), .B1(\mem[93][3] ), .B2(n7214), 
        .Z(n3168) );
  OA22D0 U4683 ( .A1(n7215), .A2(prog_data[2]), .B1(\mem[93][2] ), .B2(n7214), 
        .Z(n3167) );
  OA22D0 U4684 ( .A1(n7215), .A2(prog_data[1]), .B1(\mem[93][1] ), .B2(n7214), 
        .Z(n3166) );
  OA22D0 U4685 ( .A1(n7215), .A2(prog_data[0]), .B1(\mem[93][0] ), .B2(n7214), 
        .Z(n3165) );
  NR2D0 U4686 ( .A1(n7570), .A2(n7218), .ZN(n7216) );
  INVD0 U4687 ( .I(n7216), .ZN(n7217) );
  OA22D0 U4688 ( .A1(n7217), .A2(prog_data[15]), .B1(\mem[94][15] ), .B2(n7216), .Z(n3164) );
  OA22D0 U4689 ( .A1(n7217), .A2(prog_data[14]), .B1(\mem[94][14] ), .B2(n7216), .Z(n3163) );
  OA22D0 U4690 ( .A1(n7217), .A2(prog_data[13]), .B1(\mem[94][13] ), .B2(n7216), .Z(n3162) );
  OA22D0 U4691 ( .A1(n7217), .A2(prog_data[12]), .B1(\mem[94][12] ), .B2(n7216), .Z(n3161) );
  OA22D0 U4692 ( .A1(n7217), .A2(prog_data[11]), .B1(\mem[94][11] ), .B2(n7216), .Z(n3160) );
  OA22D0 U4693 ( .A1(n7217), .A2(prog_data[10]), .B1(\mem[94][10] ), .B2(n7216), .Z(n3159) );
  OA22D0 U4694 ( .A1(n7217), .A2(prog_data[9]), .B1(\mem[94][9] ), .B2(n7216), 
        .Z(n3158) );
  OA22D0 U4695 ( .A1(n7217), .A2(prog_data[8]), .B1(\mem[94][8] ), .B2(n7216), 
        .Z(n3157) );
  OA22D0 U4696 ( .A1(n7217), .A2(prog_data[7]), .B1(\mem[94][7] ), .B2(n7216), 
        .Z(n3156) );
  OA22D0 U4697 ( .A1(n7217), .A2(prog_data[6]), .B1(\mem[94][6] ), .B2(n7216), 
        .Z(n3155) );
  OA22D0 U4698 ( .A1(n7217), .A2(prog_data[5]), .B1(\mem[94][5] ), .B2(n7216), 
        .Z(n3154) );
  OA22D0 U4699 ( .A1(n7217), .A2(prog_data[4]), .B1(\mem[94][4] ), .B2(n7216), 
        .Z(n3153) );
  OA22D0 U4700 ( .A1(n7217), .A2(prog_data[3]), .B1(\mem[94][3] ), .B2(n7216), 
        .Z(n3152) );
  OA22D0 U4701 ( .A1(n7217), .A2(prog_data[2]), .B1(\mem[94][2] ), .B2(n7216), 
        .Z(n3151) );
  OA22D0 U4702 ( .A1(n7217), .A2(prog_data[1]), .B1(\mem[94][1] ), .B2(n7216), 
        .Z(n3150) );
  OA22D0 U4703 ( .A1(n7217), .A2(prog_data[0]), .B1(\mem[94][0] ), .B2(n7216), 
        .Z(n3149) );
  NR2D0 U4704 ( .A1(n7574), .A2(n7218), .ZN(n7219) );
  INVD0 U4705 ( .I(n7219), .ZN(n7220) );
  OA22D0 U4706 ( .A1(n7220), .A2(prog_data[15]), .B1(\mem[95][15] ), .B2(n7219), .Z(n3148) );
  OA22D0 U4707 ( .A1(n7220), .A2(prog_data[14]), .B1(\mem[95][14] ), .B2(n7219), .Z(n3147) );
  OA22D0 U4708 ( .A1(n7220), .A2(prog_data[13]), .B1(\mem[95][13] ), .B2(n7219), .Z(n3146) );
  OA22D0 U4709 ( .A1(n7220), .A2(prog_data[12]), .B1(\mem[95][12] ), .B2(n7219), .Z(n3145) );
  OA22D0 U4710 ( .A1(n7220), .A2(prog_data[11]), .B1(\mem[95][11] ), .B2(n7219), .Z(n3144) );
  OA22D0 U4711 ( .A1(n7220), .A2(prog_data[10]), .B1(\mem[95][10] ), .B2(n7219), .Z(n3143) );
  OA22D0 U4712 ( .A1(n7220), .A2(prog_data[9]), .B1(\mem[95][9] ), .B2(n7219), 
        .Z(n3142) );
  OA22D0 U4713 ( .A1(n7220), .A2(prog_data[8]), .B1(\mem[95][8] ), .B2(n7219), 
        .Z(n3141) );
  OA22D0 U4714 ( .A1(n7220), .A2(prog_data[7]), .B1(\mem[95][7] ), .B2(n7219), 
        .Z(n3140) );
  OA22D0 U4715 ( .A1(n7220), .A2(prog_data[6]), .B1(\mem[95][6] ), .B2(n7219), 
        .Z(n3139) );
  OA22D0 U4716 ( .A1(n7220), .A2(prog_data[5]), .B1(\mem[95][5] ), .B2(n7219), 
        .Z(n3138) );
  OA22D0 U4717 ( .A1(n7220), .A2(prog_data[4]), .B1(\mem[95][4] ), .B2(n7219), 
        .Z(n3137) );
  OA22D0 U4718 ( .A1(n7220), .A2(prog_data[3]), .B1(\mem[95][3] ), .B2(n7219), 
        .Z(n3136) );
  OA22D0 U4719 ( .A1(n7220), .A2(prog_data[2]), .B1(\mem[95][2] ), .B2(n7219), 
        .Z(n3135) );
  OA22D0 U4720 ( .A1(n7220), .A2(prog_data[1]), .B1(\mem[95][1] ), .B2(n7219), 
        .Z(n3134) );
  OA22D0 U4721 ( .A1(n7220), .A2(prog_data[0]), .B1(\mem[95][0] ), .B2(n7219), 
        .Z(n3133) );
  ND3D0 U4722 ( .A1(prog_addr[6]), .A2(prog_addr[5]), .A3(n7221), .ZN(n7252)
         );
  NR2D0 U4723 ( .A1(n7528), .A2(n7252), .ZN(n7222) );
  INVD0 U4724 ( .I(n7222), .ZN(n7223) );
  OA22D0 U4725 ( .A1(n7223), .A2(prog_data[15]), .B1(\mem[96][15] ), .B2(n7222), .Z(n3132) );
  OA22D0 U4726 ( .A1(n7223), .A2(prog_data[14]), .B1(\mem[96][14] ), .B2(n7222), .Z(n3131) );
  OA22D0 U4727 ( .A1(n7223), .A2(prog_data[13]), .B1(\mem[96][13] ), .B2(n7222), .Z(n3130) );
  OA22D0 U4728 ( .A1(n7223), .A2(prog_data[12]), .B1(\mem[96][12] ), .B2(n7222), .Z(n3129) );
  OA22D0 U4729 ( .A1(n7223), .A2(prog_data[11]), .B1(\mem[96][11] ), .B2(n7222), .Z(n3128) );
  OA22D0 U4730 ( .A1(n7223), .A2(prog_data[10]), .B1(\mem[96][10] ), .B2(n7222), .Z(n3127) );
  OA22D0 U4731 ( .A1(n7223), .A2(prog_data[9]), .B1(\mem[96][9] ), .B2(n7222), 
        .Z(n3126) );
  OA22D0 U4732 ( .A1(n7223), .A2(prog_data[8]), .B1(\mem[96][8] ), .B2(n7222), 
        .Z(n3125) );
  OA22D0 U4733 ( .A1(n7223), .A2(prog_data[7]), .B1(\mem[96][7] ), .B2(n7222), 
        .Z(n3124) );
  OA22D0 U4734 ( .A1(n7223), .A2(prog_data[6]), .B1(\mem[96][6] ), .B2(n7222), 
        .Z(n3123) );
  OA22D0 U4735 ( .A1(n7223), .A2(prog_data[5]), .B1(\mem[96][5] ), .B2(n7222), 
        .Z(n3122) );
  OA22D0 U4736 ( .A1(n7223), .A2(prog_data[4]), .B1(\mem[96][4] ), .B2(n7222), 
        .Z(n3121) );
  OA22D0 U4737 ( .A1(n7223), .A2(prog_data[3]), .B1(\mem[96][3] ), .B2(n7222), 
        .Z(n3120) );
  OA22D0 U4738 ( .A1(n7223), .A2(prog_data[2]), .B1(\mem[96][2] ), .B2(n7222), 
        .Z(n3119) );
  OA22D0 U4739 ( .A1(n7223), .A2(prog_data[1]), .B1(\mem[96][1] ), .B2(n7222), 
        .Z(n3118) );
  OA22D0 U4740 ( .A1(n7223), .A2(prog_data[0]), .B1(\mem[96][0] ), .B2(n7222), 
        .Z(n3117) );
  NR2D0 U4741 ( .A1(n7531), .A2(n7252), .ZN(n7224) );
  INVD0 U4742 ( .I(n7224), .ZN(n7225) );
  OA22D0 U4743 ( .A1(n7225), .A2(prog_data[15]), .B1(\mem[97][15] ), .B2(n7224), .Z(n3116) );
  OA22D0 U4744 ( .A1(n7225), .A2(prog_data[14]), .B1(\mem[97][14] ), .B2(n7224), .Z(n3115) );
  OA22D0 U4745 ( .A1(n7225), .A2(prog_data[13]), .B1(\mem[97][13] ), .B2(n7224), .Z(n3114) );
  OA22D0 U4746 ( .A1(n7225), .A2(prog_data[12]), .B1(\mem[97][12] ), .B2(n7224), .Z(n3113) );
  OA22D0 U4747 ( .A1(n7225), .A2(prog_data[11]), .B1(\mem[97][11] ), .B2(n7224), .Z(n3112) );
  OA22D0 U4748 ( .A1(n7225), .A2(prog_data[10]), .B1(\mem[97][10] ), .B2(n7224), .Z(n3111) );
  OA22D0 U4749 ( .A1(n7225), .A2(prog_data[9]), .B1(\mem[97][9] ), .B2(n7224), 
        .Z(n3110) );
  OA22D0 U4750 ( .A1(n7225), .A2(prog_data[8]), .B1(\mem[97][8] ), .B2(n7224), 
        .Z(n3109) );
  OA22D0 U4751 ( .A1(n7225), .A2(prog_data[7]), .B1(\mem[97][7] ), .B2(n7224), 
        .Z(n3108) );
  OA22D0 U4752 ( .A1(n7225), .A2(prog_data[6]), .B1(\mem[97][6] ), .B2(n7224), 
        .Z(n3107) );
  OA22D0 U4753 ( .A1(n7225), .A2(prog_data[5]), .B1(\mem[97][5] ), .B2(n7224), 
        .Z(n3106) );
  OA22D0 U4754 ( .A1(n7225), .A2(prog_data[4]), .B1(\mem[97][4] ), .B2(n7224), 
        .Z(n3105) );
  OA22D0 U4755 ( .A1(n7225), .A2(prog_data[3]), .B1(\mem[97][3] ), .B2(n7224), 
        .Z(n3104) );
  OA22D0 U4756 ( .A1(n7225), .A2(prog_data[2]), .B1(\mem[97][2] ), .B2(n7224), 
        .Z(n3103) );
  OA22D0 U4757 ( .A1(n7225), .A2(prog_data[1]), .B1(\mem[97][1] ), .B2(n7224), 
        .Z(n3102) );
  OA22D0 U4758 ( .A1(n7225), .A2(prog_data[0]), .B1(\mem[97][0] ), .B2(n7224), 
        .Z(n3101) );
  NR2D0 U4759 ( .A1(n7534), .A2(n7252), .ZN(n7226) );
  INVD0 U4760 ( .I(n7226), .ZN(n7227) );
  OA22D0 U4761 ( .A1(n7227), .A2(prog_data[15]), .B1(\mem[98][15] ), .B2(n7226), .Z(n3100) );
  OA22D0 U4762 ( .A1(n7227), .A2(prog_data[14]), .B1(\mem[98][14] ), .B2(n7226), .Z(n3099) );
  OA22D0 U4763 ( .A1(n7227), .A2(prog_data[13]), .B1(\mem[98][13] ), .B2(n7226), .Z(n3098) );
  OA22D0 U4764 ( .A1(n7227), .A2(prog_data[12]), .B1(\mem[98][12] ), .B2(n7226), .Z(n3097) );
  OA22D0 U4765 ( .A1(n7227), .A2(prog_data[11]), .B1(\mem[98][11] ), .B2(n7226), .Z(n3096) );
  OA22D0 U4766 ( .A1(n7227), .A2(prog_data[10]), .B1(\mem[98][10] ), .B2(n7226), .Z(n3095) );
  OA22D0 U4767 ( .A1(n7227), .A2(prog_data[9]), .B1(\mem[98][9] ), .B2(n7226), 
        .Z(n3094) );
  OA22D0 U4768 ( .A1(n7227), .A2(prog_data[8]), .B1(\mem[98][8] ), .B2(n7226), 
        .Z(n3093) );
  OA22D0 U4769 ( .A1(n7227), .A2(prog_data[7]), .B1(\mem[98][7] ), .B2(n7226), 
        .Z(n3092) );
  OA22D0 U4770 ( .A1(n7227), .A2(prog_data[6]), .B1(\mem[98][6] ), .B2(n7226), 
        .Z(n3091) );
  OA22D0 U4771 ( .A1(n7227), .A2(prog_data[5]), .B1(\mem[98][5] ), .B2(n7226), 
        .Z(n3090) );
  OA22D0 U4772 ( .A1(n7227), .A2(prog_data[4]), .B1(\mem[98][4] ), .B2(n7226), 
        .Z(n3089) );
  OA22D0 U4773 ( .A1(n7227), .A2(prog_data[3]), .B1(\mem[98][3] ), .B2(n7226), 
        .Z(n3088) );
  OA22D0 U4774 ( .A1(n7227), .A2(prog_data[2]), .B1(\mem[98][2] ), .B2(n7226), 
        .Z(n3087) );
  OA22D0 U4775 ( .A1(n7227), .A2(prog_data[1]), .B1(\mem[98][1] ), .B2(n7226), 
        .Z(n3086) );
  OA22D0 U4776 ( .A1(n7227), .A2(prog_data[0]), .B1(\mem[98][0] ), .B2(n7226), 
        .Z(n3085) );
  NR2D0 U4777 ( .A1(n7537), .A2(n7252), .ZN(n7228) );
  OA22D0 U4778 ( .A1(n7229), .A2(prog_data[15]), .B1(\mem[99][15] ), .B2(n7228), .Z(n3084) );
  OA22D0 U4779 ( .A1(n7229), .A2(prog_data[14]), .B1(\mem[99][14] ), .B2(n7228), .Z(n3083) );
  OA22D0 U4780 ( .A1(n7229), .A2(prog_data[13]), .B1(\mem[99][13] ), .B2(n7228), .Z(n3082) );
  OA22D0 U4781 ( .A1(n7229), .A2(prog_data[12]), .B1(\mem[99][12] ), .B2(n7228), .Z(n3081) );
  OA22D0 U4782 ( .A1(n7229), .A2(prog_data[11]), .B1(\mem[99][11] ), .B2(n7228), .Z(n3080) );
  OA22D0 U4783 ( .A1(n7229), .A2(prog_data[10]), .B1(\mem[99][10] ), .B2(n7228), .Z(n3079) );
  OA22D0 U4784 ( .A1(n7229), .A2(prog_data[9]), .B1(\mem[99][9] ), .B2(n7228), 
        .Z(n3078) );
  OA22D0 U4785 ( .A1(n7229), .A2(prog_data[8]), .B1(\mem[99][8] ), .B2(n7228), 
        .Z(n3077) );
  OA22D0 U4786 ( .A1(n7229), .A2(prog_data[7]), .B1(\mem[99][7] ), .B2(n7228), 
        .Z(n3076) );
  OA22D0 U4787 ( .A1(n7229), .A2(prog_data[6]), .B1(\mem[99][6] ), .B2(n7228), 
        .Z(n3075) );
  OA22D0 U4788 ( .A1(n7229), .A2(prog_data[5]), .B1(\mem[99][5] ), .B2(n7228), 
        .Z(n3074) );
  OA22D0 U4789 ( .A1(n7229), .A2(prog_data[4]), .B1(\mem[99][4] ), .B2(n7228), 
        .Z(n3073) );
  OA22D0 U4790 ( .A1(n7229), .A2(prog_data[3]), .B1(\mem[99][3] ), .B2(n7228), 
        .Z(n3072) );
  OA22D0 U4791 ( .A1(n7229), .A2(prog_data[2]), .B1(\mem[99][2] ), .B2(n7228), 
        .Z(n3071) );
  OA22D0 U4792 ( .A1(n7229), .A2(prog_data[1]), .B1(\mem[99][1] ), .B2(n7228), 
        .Z(n3070) );
  OA22D0 U4793 ( .A1(n7229), .A2(prog_data[0]), .B1(\mem[99][0] ), .B2(n7228), 
        .Z(n3069) );
  NR2D0 U4794 ( .A1(n7540), .A2(n7252), .ZN(n7230) );
  INVD0 U4795 ( .I(n7230), .ZN(n7231) );
  OA22D0 U4796 ( .A1(n7231), .A2(prog_data[15]), .B1(\mem[100][15] ), .B2(
        n7230), .Z(n3068) );
  OA22D0 U4797 ( .A1(n7231), .A2(prog_data[14]), .B1(\mem[100][14] ), .B2(
        n7230), .Z(n3067) );
  OA22D0 U4798 ( .A1(n7231), .A2(prog_data[13]), .B1(\mem[100][13] ), .B2(
        n7230), .Z(n3066) );
  OA22D0 U4799 ( .A1(n7231), .A2(prog_data[12]), .B1(\mem[100][12] ), .B2(
        n7230), .Z(n3065) );
  OA22D0 U4800 ( .A1(n7231), .A2(prog_data[11]), .B1(\mem[100][11] ), .B2(
        n7230), .Z(n3064) );
  OA22D0 U4801 ( .A1(n7231), .A2(prog_data[10]), .B1(\mem[100][10] ), .B2(
        n7230), .Z(n3063) );
  OA22D0 U4802 ( .A1(n7231), .A2(prog_data[9]), .B1(\mem[100][9] ), .B2(n7230), 
        .Z(n3062) );
  OA22D0 U4803 ( .A1(n7231), .A2(prog_data[8]), .B1(\mem[100][8] ), .B2(n7230), 
        .Z(n3061) );
  OA22D0 U4804 ( .A1(n7231), .A2(prog_data[7]), .B1(\mem[100][7] ), .B2(n7230), 
        .Z(n3060) );
  OA22D0 U4805 ( .A1(n7231), .A2(prog_data[6]), .B1(\mem[100][6] ), .B2(n7230), 
        .Z(n3059) );
  OA22D0 U4806 ( .A1(n7231), .A2(prog_data[5]), .B1(\mem[100][5] ), .B2(n7230), 
        .Z(n3058) );
  OA22D0 U4807 ( .A1(n7231), .A2(prog_data[4]), .B1(\mem[100][4] ), .B2(n7230), 
        .Z(n3057) );
  OA22D0 U4808 ( .A1(n7231), .A2(prog_data[3]), .B1(\mem[100][3] ), .B2(n7230), 
        .Z(n3056) );
  OA22D0 U4809 ( .A1(n7231), .A2(prog_data[2]), .B1(\mem[100][2] ), .B2(n7230), 
        .Z(n3055) );
  OA22D0 U4810 ( .A1(n7231), .A2(prog_data[1]), .B1(\mem[100][1] ), .B2(n7230), 
        .Z(n3054) );
  OA22D0 U4811 ( .A1(n7231), .A2(prog_data[0]), .B1(\mem[100][0] ), .B2(n7230), 
        .Z(n3053) );
  NR2D0 U4812 ( .A1(n7543), .A2(n7252), .ZN(n7232) );
  INVD0 U4813 ( .I(n7232), .ZN(n7233) );
  OA22D0 U4814 ( .A1(n7233), .A2(prog_data[15]), .B1(\mem[101][15] ), .B2(
        n7232), .Z(n3052) );
  OA22D0 U4815 ( .A1(n7233), .A2(prog_data[14]), .B1(\mem[101][14] ), .B2(
        n7232), .Z(n3051) );
  OA22D0 U4816 ( .A1(n7233), .A2(prog_data[13]), .B1(\mem[101][13] ), .B2(
        n7232), .Z(n3050) );
  OA22D0 U4817 ( .A1(n7233), .A2(prog_data[12]), .B1(\mem[101][12] ), .B2(
        n7232), .Z(n3049) );
  OA22D0 U4818 ( .A1(n7233), .A2(prog_data[11]), .B1(\mem[101][11] ), .B2(
        n7232), .Z(n3048) );
  OA22D0 U4819 ( .A1(n7233), .A2(prog_data[10]), .B1(\mem[101][10] ), .B2(
        n7232), .Z(n3047) );
  OA22D0 U4820 ( .A1(n7233), .A2(prog_data[9]), .B1(\mem[101][9] ), .B2(n7232), 
        .Z(n3046) );
  OA22D0 U4821 ( .A1(n7233), .A2(prog_data[8]), .B1(\mem[101][8] ), .B2(n7232), 
        .Z(n3045) );
  OA22D0 U4822 ( .A1(n7233), .A2(prog_data[7]), .B1(\mem[101][7] ), .B2(n7232), 
        .Z(n3044) );
  OA22D0 U4823 ( .A1(n7233), .A2(prog_data[6]), .B1(\mem[101][6] ), .B2(n7232), 
        .Z(n3043) );
  OA22D0 U4824 ( .A1(n7233), .A2(prog_data[5]), .B1(\mem[101][5] ), .B2(n7232), 
        .Z(n3042) );
  OA22D0 U4825 ( .A1(n7233), .A2(prog_data[4]), .B1(\mem[101][4] ), .B2(n7232), 
        .Z(n3041) );
  OA22D0 U4826 ( .A1(n7233), .A2(prog_data[3]), .B1(\mem[101][3] ), .B2(n7232), 
        .Z(n3040) );
  OA22D0 U4827 ( .A1(n7233), .A2(prog_data[2]), .B1(\mem[101][2] ), .B2(n7232), 
        .Z(n3039) );
  OA22D0 U4828 ( .A1(n7233), .A2(prog_data[1]), .B1(\mem[101][1] ), .B2(n7232), 
        .Z(n3038) );
  OA22D0 U4829 ( .A1(n7233), .A2(prog_data[0]), .B1(\mem[101][0] ), .B2(n7232), 
        .Z(n3037) );
  NR2D0 U4830 ( .A1(n7546), .A2(n7252), .ZN(n7234) );
  INVD0 U4831 ( .I(n7234), .ZN(n7235) );
  OA22D0 U4832 ( .A1(n7235), .A2(prog_data[15]), .B1(\mem[102][15] ), .B2(
        n7234), .Z(n3036) );
  OA22D0 U4833 ( .A1(n7235), .A2(prog_data[14]), .B1(\mem[102][14] ), .B2(
        n7234), .Z(n3035) );
  OA22D0 U4834 ( .A1(n7235), .A2(prog_data[13]), .B1(\mem[102][13] ), .B2(
        n7234), .Z(n3034) );
  OA22D0 U4835 ( .A1(n7235), .A2(prog_data[12]), .B1(\mem[102][12] ), .B2(
        n7234), .Z(n3033) );
  OA22D0 U4836 ( .A1(n7235), .A2(prog_data[11]), .B1(\mem[102][11] ), .B2(
        n7234), .Z(n3032) );
  OA22D0 U4837 ( .A1(n7235), .A2(prog_data[10]), .B1(\mem[102][10] ), .B2(
        n7234), .Z(n3031) );
  OA22D0 U4838 ( .A1(n7235), .A2(prog_data[9]), .B1(\mem[102][9] ), .B2(n7234), 
        .Z(n3030) );
  OA22D0 U4839 ( .A1(n7235), .A2(prog_data[8]), .B1(\mem[102][8] ), .B2(n7234), 
        .Z(n3029) );
  OA22D0 U4840 ( .A1(n7235), .A2(prog_data[7]), .B1(\mem[102][7] ), .B2(n7234), 
        .Z(n3028) );
  OA22D0 U4841 ( .A1(n7235), .A2(prog_data[6]), .B1(\mem[102][6] ), .B2(n7234), 
        .Z(n3027) );
  OA22D0 U4842 ( .A1(n7235), .A2(prog_data[5]), .B1(\mem[102][5] ), .B2(n7234), 
        .Z(n3026) );
  OA22D0 U4843 ( .A1(n7235), .A2(prog_data[4]), .B1(\mem[102][4] ), .B2(n7234), 
        .Z(n3025) );
  OA22D0 U4844 ( .A1(n7235), .A2(prog_data[3]), .B1(\mem[102][3] ), .B2(n7234), 
        .Z(n3024) );
  OA22D0 U4845 ( .A1(n7235), .A2(prog_data[2]), .B1(\mem[102][2] ), .B2(n7234), 
        .Z(n3023) );
  OA22D0 U4846 ( .A1(n7235), .A2(prog_data[1]), .B1(\mem[102][1] ), .B2(n7234), 
        .Z(n3022) );
  OA22D0 U4847 ( .A1(n7235), .A2(prog_data[0]), .B1(\mem[102][0] ), .B2(n7234), 
        .Z(n3021) );
  NR2D0 U4848 ( .A1(n7549), .A2(n7252), .ZN(n7236) );
  INVD0 U4849 ( .I(n7236), .ZN(n7237) );
  OA22D0 U4850 ( .A1(n7237), .A2(prog_data[15]), .B1(\mem[103][15] ), .B2(
        n7236), .Z(n3020) );
  OA22D0 U4851 ( .A1(n7237), .A2(prog_data[14]), .B1(\mem[103][14] ), .B2(
        n7236), .Z(n3019) );
  OA22D0 U4852 ( .A1(n7237), .A2(prog_data[13]), .B1(\mem[103][13] ), .B2(
        n7236), .Z(n3018) );
  OA22D0 U4853 ( .A1(n7237), .A2(prog_data[12]), .B1(\mem[103][12] ), .B2(
        n7236), .Z(n3017) );
  OA22D0 U4854 ( .A1(n7237), .A2(prog_data[11]), .B1(\mem[103][11] ), .B2(
        n7236), .Z(n3016) );
  OA22D0 U4855 ( .A1(n7237), .A2(prog_data[10]), .B1(\mem[103][10] ), .B2(
        n7236), .Z(n3015) );
  OA22D0 U4856 ( .A1(n7237), .A2(prog_data[9]), .B1(\mem[103][9] ), .B2(n7236), 
        .Z(n3014) );
  OA22D0 U4857 ( .A1(n7237), .A2(prog_data[8]), .B1(\mem[103][8] ), .B2(n7236), 
        .Z(n3013) );
  OA22D0 U4858 ( .A1(n7237), .A2(prog_data[7]), .B1(\mem[103][7] ), .B2(n7236), 
        .Z(n3012) );
  OA22D0 U4859 ( .A1(n7237), .A2(prog_data[6]), .B1(\mem[103][6] ), .B2(n7236), 
        .Z(n3011) );
  OA22D0 U4860 ( .A1(n7237), .A2(prog_data[5]), .B1(\mem[103][5] ), .B2(n7236), 
        .Z(n3010) );
  OA22D0 U4861 ( .A1(n7237), .A2(prog_data[4]), .B1(\mem[103][4] ), .B2(n7236), 
        .Z(n3009) );
  OA22D0 U4862 ( .A1(n7237), .A2(prog_data[3]), .B1(\mem[103][3] ), .B2(n7236), 
        .Z(n3008) );
  OA22D0 U4863 ( .A1(n7237), .A2(prog_data[2]), .B1(\mem[103][2] ), .B2(n7236), 
        .Z(n3007) );
  OA22D0 U4864 ( .A1(n7237), .A2(prog_data[1]), .B1(\mem[103][1] ), .B2(n7236), 
        .Z(n3006) );
  OA22D0 U4865 ( .A1(n7237), .A2(prog_data[0]), .B1(\mem[103][0] ), .B2(n7236), 
        .Z(n3005) );
  NR2D0 U4866 ( .A1(n7552), .A2(n7252), .ZN(n7238) );
  INVD0 U4867 ( .I(n7238), .ZN(n7239) );
  OA22D0 U4868 ( .A1(n7239), .A2(prog_data[15]), .B1(\mem[104][15] ), .B2(
        n7238), .Z(n3004) );
  OA22D0 U4869 ( .A1(n7239), .A2(prog_data[14]), .B1(\mem[104][14] ), .B2(
        n7238), .Z(n3003) );
  OA22D0 U4870 ( .A1(n7239), .A2(prog_data[13]), .B1(\mem[104][13] ), .B2(
        n7238), .Z(n3002) );
  OA22D0 U4871 ( .A1(n7239), .A2(prog_data[12]), .B1(\mem[104][12] ), .B2(
        n7238), .Z(n3001) );
  OA22D0 U4872 ( .A1(n7239), .A2(prog_data[11]), .B1(\mem[104][11] ), .B2(
        n7238), .Z(n3000) );
  OA22D0 U4873 ( .A1(n7239), .A2(prog_data[10]), .B1(\mem[104][10] ), .B2(
        n7238), .Z(n2999) );
  OA22D0 U4874 ( .A1(n7239), .A2(prog_data[9]), .B1(\mem[104][9] ), .B2(n7238), 
        .Z(n2998) );
  OA22D0 U4875 ( .A1(n7239), .A2(prog_data[8]), .B1(\mem[104][8] ), .B2(n7238), 
        .Z(n2997) );
  OA22D0 U4876 ( .A1(n7239), .A2(prog_data[7]), .B1(\mem[104][7] ), .B2(n7238), 
        .Z(n2996) );
  OA22D0 U4877 ( .A1(n7239), .A2(prog_data[6]), .B1(\mem[104][6] ), .B2(n7238), 
        .Z(n2995) );
  OA22D0 U4878 ( .A1(n7239), .A2(prog_data[5]), .B1(\mem[104][5] ), .B2(n7238), 
        .Z(n2994) );
  OA22D0 U4879 ( .A1(n7239), .A2(prog_data[4]), .B1(\mem[104][4] ), .B2(n7238), 
        .Z(n2993) );
  OA22D0 U4880 ( .A1(n7239), .A2(prog_data[3]), .B1(\mem[104][3] ), .B2(n7238), 
        .Z(n2992) );
  OA22D0 U4881 ( .A1(n7239), .A2(prog_data[2]), .B1(\mem[104][2] ), .B2(n7238), 
        .Z(n2991) );
  OA22D0 U4882 ( .A1(n7239), .A2(prog_data[1]), .B1(\mem[104][1] ), .B2(n7238), 
        .Z(n2990) );
  OA22D0 U4883 ( .A1(n7239), .A2(prog_data[0]), .B1(\mem[104][0] ), .B2(n7238), 
        .Z(n2989) );
  NR2D0 U4884 ( .A1(n7555), .A2(n7252), .ZN(n7240) );
  INVD0 U4885 ( .I(n7240), .ZN(n7241) );
  OA22D0 U4886 ( .A1(n7241), .A2(prog_data[15]), .B1(\mem[105][15] ), .B2(
        n7240), .Z(n2988) );
  OA22D0 U4887 ( .A1(n7241), .A2(prog_data[14]), .B1(\mem[105][14] ), .B2(
        n7240), .Z(n2987) );
  OA22D0 U4888 ( .A1(n7241), .A2(prog_data[13]), .B1(\mem[105][13] ), .B2(
        n7240), .Z(n2986) );
  OA22D0 U4889 ( .A1(n7241), .A2(prog_data[12]), .B1(\mem[105][12] ), .B2(
        n7240), .Z(n2985) );
  OA22D0 U4890 ( .A1(n7241), .A2(prog_data[11]), .B1(\mem[105][11] ), .B2(
        n7240), .Z(n2984) );
  OA22D0 U4891 ( .A1(n7241), .A2(prog_data[10]), .B1(\mem[105][10] ), .B2(
        n7240), .Z(n2983) );
  OA22D0 U4892 ( .A1(n7241), .A2(prog_data[9]), .B1(\mem[105][9] ), .B2(n7240), 
        .Z(n2982) );
  OA22D0 U4893 ( .A1(n7241), .A2(prog_data[8]), .B1(\mem[105][8] ), .B2(n7240), 
        .Z(n2981) );
  OA22D0 U4894 ( .A1(n7241), .A2(prog_data[7]), .B1(\mem[105][7] ), .B2(n7240), 
        .Z(n2980) );
  OA22D0 U4895 ( .A1(n7241), .A2(prog_data[6]), .B1(\mem[105][6] ), .B2(n7240), 
        .Z(n2979) );
  OA22D0 U4896 ( .A1(n7241), .A2(prog_data[5]), .B1(\mem[105][5] ), .B2(n7240), 
        .Z(n2978) );
  OA22D0 U4897 ( .A1(n7241), .A2(prog_data[4]), .B1(\mem[105][4] ), .B2(n7240), 
        .Z(n2977) );
  OA22D0 U4898 ( .A1(n7241), .A2(prog_data[3]), .B1(\mem[105][3] ), .B2(n7240), 
        .Z(n2976) );
  OA22D0 U4899 ( .A1(n7241), .A2(prog_data[2]), .B1(\mem[105][2] ), .B2(n7240), 
        .Z(n2975) );
  OA22D0 U4900 ( .A1(n7241), .A2(prog_data[1]), .B1(\mem[105][1] ), .B2(n7240), 
        .Z(n2974) );
  OA22D0 U4901 ( .A1(n7241), .A2(prog_data[0]), .B1(\mem[105][0] ), .B2(n7240), 
        .Z(n2973) );
  INVD0 U4902 ( .I(n7242), .ZN(n7243) );
  OA22D0 U4903 ( .A1(n7243), .A2(prog_data[15]), .B1(\mem[106][15] ), .B2(
        n7242), .Z(n2972) );
  OA22D0 U4904 ( .A1(n7243), .A2(prog_data[14]), .B1(\mem[106][14] ), .B2(
        n7242), .Z(n2971) );
  OA22D0 U4905 ( .A1(n7243), .A2(prog_data[13]), .B1(\mem[106][13] ), .B2(
        n7242), .Z(n2970) );
  OA22D0 U4906 ( .A1(n7243), .A2(prog_data[12]), .B1(\mem[106][12] ), .B2(
        n7242), .Z(n2969) );
  OA22D0 U4907 ( .A1(n7243), .A2(prog_data[11]), .B1(\mem[106][11] ), .B2(
        n7242), .Z(n2968) );
  OA22D0 U4908 ( .A1(n7243), .A2(prog_data[10]), .B1(\mem[106][10] ), .B2(
        n7242), .Z(n2967) );
  OA22D0 U4909 ( .A1(n7243), .A2(prog_data[9]), .B1(\mem[106][9] ), .B2(n7242), 
        .Z(n2966) );
  OA22D0 U4910 ( .A1(n7243), .A2(prog_data[8]), .B1(\mem[106][8] ), .B2(n7242), 
        .Z(n2965) );
  OA22D0 U4911 ( .A1(n7243), .A2(prog_data[7]), .B1(\mem[106][7] ), .B2(n7242), 
        .Z(n2964) );
  OA22D0 U4912 ( .A1(n7243), .A2(prog_data[6]), .B1(\mem[106][6] ), .B2(n7242), 
        .Z(n2963) );
  OA22D0 U4913 ( .A1(n7243), .A2(prog_data[5]), .B1(\mem[106][5] ), .B2(n7242), 
        .Z(n2962) );
  OA22D0 U4914 ( .A1(n7243), .A2(prog_data[4]), .B1(\mem[106][4] ), .B2(n7242), 
        .Z(n2961) );
  OA22D0 U4915 ( .A1(n7243), .A2(prog_data[3]), .B1(\mem[106][3] ), .B2(n7242), 
        .Z(n2960) );
  OA22D0 U4916 ( .A1(n7243), .A2(prog_data[2]), .B1(\mem[106][2] ), .B2(n7242), 
        .Z(n2959) );
  OA22D0 U4917 ( .A1(n7243), .A2(prog_data[1]), .B1(\mem[106][1] ), .B2(n7242), 
        .Z(n2958) );
  OA22D0 U4918 ( .A1(n7243), .A2(prog_data[0]), .B1(\mem[106][0] ), .B2(n7242), 
        .Z(n2957) );
  NR2D0 U4919 ( .A1(n7561), .A2(n7252), .ZN(n7244) );
  INVD0 U4920 ( .I(n7244), .ZN(n7245) );
  OA22D0 U4921 ( .A1(n7245), .A2(prog_data[15]), .B1(\mem[107][15] ), .B2(
        n7244), .Z(n2956) );
  OA22D0 U4922 ( .A1(n7245), .A2(prog_data[14]), .B1(\mem[107][14] ), .B2(
        n7244), .Z(n2955) );
  OA22D0 U4923 ( .A1(n7245), .A2(prog_data[13]), .B1(\mem[107][13] ), .B2(
        n7244), .Z(n2954) );
  OA22D0 U4924 ( .A1(n7245), .A2(prog_data[12]), .B1(\mem[107][12] ), .B2(
        n7244), .Z(n2953) );
  OA22D0 U4925 ( .A1(n7245), .A2(prog_data[11]), .B1(\mem[107][11] ), .B2(
        n7244), .Z(n2952) );
  OA22D0 U4926 ( .A1(n7245), .A2(prog_data[10]), .B1(\mem[107][10] ), .B2(
        n7244), .Z(n2951) );
  OA22D0 U4927 ( .A1(n7245), .A2(prog_data[9]), .B1(\mem[107][9] ), .B2(n7244), 
        .Z(n2950) );
  OA22D0 U4928 ( .A1(n7245), .A2(prog_data[8]), .B1(\mem[107][8] ), .B2(n7244), 
        .Z(n2949) );
  OA22D0 U4929 ( .A1(n7245), .A2(prog_data[7]), .B1(\mem[107][7] ), .B2(n7244), 
        .Z(n2948) );
  OA22D0 U4930 ( .A1(n7245), .A2(prog_data[6]), .B1(\mem[107][6] ), .B2(n7244), 
        .Z(n2947) );
  OA22D0 U4931 ( .A1(n7245), .A2(prog_data[5]), .B1(\mem[107][5] ), .B2(n7244), 
        .Z(n2946) );
  OA22D0 U4932 ( .A1(n7245), .A2(prog_data[4]), .B1(\mem[107][4] ), .B2(n7244), 
        .Z(n2945) );
  OA22D0 U4933 ( .A1(n7245), .A2(prog_data[3]), .B1(\mem[107][3] ), .B2(n7244), 
        .Z(n2944) );
  OA22D0 U4934 ( .A1(n7245), .A2(prog_data[2]), .B1(\mem[107][2] ), .B2(n7244), 
        .Z(n2943) );
  OA22D0 U4935 ( .A1(n7245), .A2(prog_data[1]), .B1(\mem[107][1] ), .B2(n7244), 
        .Z(n2942) );
  OA22D0 U4936 ( .A1(n7245), .A2(prog_data[0]), .B1(\mem[107][0] ), .B2(n7244), 
        .Z(n2941) );
  NR2D0 U4937 ( .A1(n7564), .A2(n7252), .ZN(n7246) );
  INVD0 U4938 ( .I(n7246), .ZN(n7247) );
  OA22D0 U4939 ( .A1(n7247), .A2(prog_data[15]), .B1(\mem[108][15] ), .B2(
        n7246), .Z(n2940) );
  OA22D0 U4940 ( .A1(n7247), .A2(prog_data[14]), .B1(\mem[108][14] ), .B2(
        n7246), .Z(n2939) );
  OA22D0 U4941 ( .A1(n7247), .A2(prog_data[13]), .B1(\mem[108][13] ), .B2(
        n7246), .Z(n2938) );
  OA22D0 U4942 ( .A1(n7247), .A2(prog_data[12]), .B1(\mem[108][12] ), .B2(
        n7246), .Z(n2937) );
  OA22D0 U4943 ( .A1(n7247), .A2(prog_data[11]), .B1(\mem[108][11] ), .B2(
        n7246), .Z(n2936) );
  OA22D0 U4944 ( .A1(n7247), .A2(prog_data[10]), .B1(\mem[108][10] ), .B2(
        n7246), .Z(n2935) );
  OA22D0 U4945 ( .A1(n7247), .A2(prog_data[9]), .B1(\mem[108][9] ), .B2(n7246), 
        .Z(n2934) );
  OA22D0 U4946 ( .A1(n7247), .A2(prog_data[8]), .B1(\mem[108][8] ), .B2(n7246), 
        .Z(n2933) );
  OA22D0 U4947 ( .A1(n7247), .A2(prog_data[7]), .B1(\mem[108][7] ), .B2(n7246), 
        .Z(n2932) );
  OA22D0 U4948 ( .A1(n7247), .A2(prog_data[6]), .B1(\mem[108][6] ), .B2(n7246), 
        .Z(n2931) );
  OA22D0 U4949 ( .A1(n7247), .A2(prog_data[5]), .B1(\mem[108][5] ), .B2(n7246), 
        .Z(n2930) );
  OA22D0 U4950 ( .A1(n7247), .A2(prog_data[4]), .B1(\mem[108][4] ), .B2(n7246), 
        .Z(n2929) );
  OA22D0 U4951 ( .A1(n7247), .A2(prog_data[3]), .B1(\mem[108][3] ), .B2(n7246), 
        .Z(n2928) );
  OA22D0 U4952 ( .A1(n7247), .A2(prog_data[2]), .B1(\mem[108][2] ), .B2(n7246), 
        .Z(n2927) );
  OA22D0 U4953 ( .A1(n7247), .A2(prog_data[1]), .B1(\mem[108][1] ), .B2(n7246), 
        .Z(n2926) );
  OA22D0 U4954 ( .A1(n7247), .A2(prog_data[0]), .B1(\mem[108][0] ), .B2(n7246), 
        .Z(n2925) );
  NR2D0 U4955 ( .A1(n7567), .A2(n7252), .ZN(n7248) );
  INVD0 U4956 ( .I(n7248), .ZN(n7249) );
  OA22D0 U4957 ( .A1(n7249), .A2(prog_data[15]), .B1(\mem[109][15] ), .B2(
        n7248), .Z(n2924) );
  OA22D0 U4958 ( .A1(n7249), .A2(prog_data[14]), .B1(\mem[109][14] ), .B2(
        n7248), .Z(n2923) );
  OA22D0 U4959 ( .A1(n7249), .A2(prog_data[13]), .B1(\mem[109][13] ), .B2(
        n7248), .Z(n2922) );
  OA22D0 U4960 ( .A1(n7249), .A2(prog_data[12]), .B1(\mem[109][12] ), .B2(
        n7248), .Z(n2921) );
  OA22D0 U4961 ( .A1(n7249), .A2(prog_data[11]), .B1(\mem[109][11] ), .B2(
        n7248), .Z(n2920) );
  OA22D0 U4962 ( .A1(n7249), .A2(prog_data[10]), .B1(\mem[109][10] ), .B2(
        n7248), .Z(n2919) );
  OA22D0 U4963 ( .A1(n7249), .A2(prog_data[9]), .B1(\mem[109][9] ), .B2(n7248), 
        .Z(n2918) );
  OA22D0 U4964 ( .A1(n7249), .A2(prog_data[8]), .B1(\mem[109][8] ), .B2(n7248), 
        .Z(n2917) );
  OA22D0 U4965 ( .A1(n7249), .A2(prog_data[7]), .B1(\mem[109][7] ), .B2(n7248), 
        .Z(n2916) );
  OA22D0 U4966 ( .A1(n7249), .A2(prog_data[6]), .B1(\mem[109][6] ), .B2(n7248), 
        .Z(n2915) );
  OA22D0 U4967 ( .A1(n7249), .A2(prog_data[5]), .B1(\mem[109][5] ), .B2(n7248), 
        .Z(n2914) );
  OA22D0 U4968 ( .A1(n7249), .A2(prog_data[4]), .B1(\mem[109][4] ), .B2(n7248), 
        .Z(n2913) );
  OA22D0 U4969 ( .A1(n7249), .A2(prog_data[3]), .B1(\mem[109][3] ), .B2(n7248), 
        .Z(n2912) );
  OA22D0 U4970 ( .A1(n7249), .A2(prog_data[2]), .B1(\mem[109][2] ), .B2(n7248), 
        .Z(n2911) );
  OA22D0 U4971 ( .A1(n7249), .A2(prog_data[1]), .B1(\mem[109][1] ), .B2(n7248), 
        .Z(n2910) );
  OA22D0 U4972 ( .A1(n7249), .A2(prog_data[0]), .B1(\mem[109][0] ), .B2(n7248), 
        .Z(n2909) );
  NR2D0 U4973 ( .A1(n7570), .A2(n7252), .ZN(n7250) );
  INVD0 U4974 ( .I(n7250), .ZN(n7251) );
  OA22D0 U4975 ( .A1(n7251), .A2(prog_data[15]), .B1(\mem[110][15] ), .B2(
        n7250), .Z(n2908) );
  OA22D0 U4976 ( .A1(n7251), .A2(prog_data[14]), .B1(\mem[110][14] ), .B2(
        n7250), .Z(n2907) );
  OA22D0 U4977 ( .A1(n7251), .A2(prog_data[13]), .B1(\mem[110][13] ), .B2(
        n7250), .Z(n2906) );
  OA22D0 U4978 ( .A1(n7251), .A2(prog_data[12]), .B1(\mem[110][12] ), .B2(
        n7250), .Z(n2905) );
  OA22D0 U4979 ( .A1(n7251), .A2(prog_data[11]), .B1(\mem[110][11] ), .B2(
        n7250), .Z(n2904) );
  OA22D0 U4980 ( .A1(n7251), .A2(prog_data[10]), .B1(\mem[110][10] ), .B2(
        n7250), .Z(n2903) );
  OA22D0 U4981 ( .A1(n7251), .A2(prog_data[9]), .B1(\mem[110][9] ), .B2(n7250), 
        .Z(n2902) );
  OA22D0 U4982 ( .A1(n7251), .A2(prog_data[8]), .B1(\mem[110][8] ), .B2(n7250), 
        .Z(n2901) );
  OA22D0 U4983 ( .A1(n7251), .A2(prog_data[7]), .B1(\mem[110][7] ), .B2(n7250), 
        .Z(n2900) );
  OA22D0 U4984 ( .A1(n7251), .A2(prog_data[6]), .B1(\mem[110][6] ), .B2(n7250), 
        .Z(n2899) );
  OA22D0 U4985 ( .A1(n7251), .A2(prog_data[5]), .B1(\mem[110][5] ), .B2(n7250), 
        .Z(n2898) );
  OA22D0 U4986 ( .A1(n7251), .A2(prog_data[4]), .B1(\mem[110][4] ), .B2(n7250), 
        .Z(n2897) );
  OA22D0 U4987 ( .A1(n7251), .A2(prog_data[3]), .B1(\mem[110][3] ), .B2(n7250), 
        .Z(n2896) );
  OA22D0 U4988 ( .A1(n7251), .A2(prog_data[2]), .B1(\mem[110][2] ), .B2(n7250), 
        .Z(n2895) );
  OA22D0 U4989 ( .A1(n7251), .A2(prog_data[1]), .B1(\mem[110][1] ), .B2(n7250), 
        .Z(n2894) );
  OA22D0 U4990 ( .A1(n7251), .A2(prog_data[0]), .B1(\mem[110][0] ), .B2(n7250), 
        .Z(n2893) );
  NR2D0 U4991 ( .A1(n7574), .A2(n7252), .ZN(n7253) );
  INVD0 U4992 ( .I(n7253), .ZN(n7254) );
  OA22D0 U4993 ( .A1(n7254), .A2(prog_data[15]), .B1(\mem[111][15] ), .B2(
        n7253), .Z(n2892) );
  OA22D0 U4994 ( .A1(n7254), .A2(prog_data[14]), .B1(\mem[111][14] ), .B2(
        n7253), .Z(n2891) );
  OA22D0 U4995 ( .A1(n7254), .A2(prog_data[13]), .B1(\mem[111][13] ), .B2(
        n7253), .Z(n2890) );
  OA22D0 U4996 ( .A1(n7254), .A2(prog_data[12]), .B1(\mem[111][12] ), .B2(
        n7253), .Z(n2889) );
  OA22D0 U4997 ( .A1(n7254), .A2(prog_data[11]), .B1(\mem[111][11] ), .B2(
        n7253), .Z(n2888) );
  OA22D0 U4998 ( .A1(n7254), .A2(prog_data[10]), .B1(\mem[111][10] ), .B2(
        n7253), .Z(n2887) );
  OA22D0 U4999 ( .A1(n7254), .A2(prog_data[9]), .B1(\mem[111][9] ), .B2(n7253), 
        .Z(n2886) );
  OA22D0 U5000 ( .A1(n7254), .A2(prog_data[8]), .B1(\mem[111][8] ), .B2(n7253), 
        .Z(n2885) );
  OA22D0 U5001 ( .A1(n7254), .A2(prog_data[7]), .B1(\mem[111][7] ), .B2(n7253), 
        .Z(n2884) );
  OA22D0 U5002 ( .A1(n7254), .A2(prog_data[6]), .B1(\mem[111][6] ), .B2(n7253), 
        .Z(n2883) );
  OA22D0 U5003 ( .A1(n7254), .A2(prog_data[5]), .B1(\mem[111][5] ), .B2(n7253), 
        .Z(n2882) );
  OA22D0 U5004 ( .A1(n7254), .A2(prog_data[4]), .B1(\mem[111][4] ), .B2(n7253), 
        .Z(n2881) );
  OA22D0 U5005 ( .A1(n7254), .A2(prog_data[3]), .B1(\mem[111][3] ), .B2(n7253), 
        .Z(n2880) );
  OA22D0 U5006 ( .A1(n7254), .A2(prog_data[2]), .B1(\mem[111][2] ), .B2(n7253), 
        .Z(n2879) );
  OA22D0 U5007 ( .A1(n7254), .A2(prog_data[1]), .B1(\mem[111][1] ), .B2(n7253), 
        .Z(n2878) );
  OA22D0 U5008 ( .A1(n7254), .A2(prog_data[0]), .B1(\mem[111][0] ), .B2(n7253), 
        .Z(n2877) );
  ND3D0 U5009 ( .A1(prog_addr[6]), .A2(prog_addr[5]), .A3(n7255), .ZN(n7286)
         );
  NR2D0 U5010 ( .A1(n7528), .A2(n7286), .ZN(n7256) );
  INVD0 U5011 ( .I(n7256), .ZN(n7257) );
  OA22D0 U5012 ( .A1(n7257), .A2(prog_data[15]), .B1(\mem[112][15] ), .B2(
        n7256), .Z(n2876) );
  OA22D0 U5013 ( .A1(n7257), .A2(prog_data[14]), .B1(\mem[112][14] ), .B2(
        n7256), .Z(n2875) );
  OA22D0 U5014 ( .A1(n7257), .A2(prog_data[13]), .B1(\mem[112][13] ), .B2(
        n7256), .Z(n2874) );
  OA22D0 U5015 ( .A1(n7257), .A2(prog_data[12]), .B1(\mem[112][12] ), .B2(
        n7256), .Z(n2873) );
  OA22D0 U5016 ( .A1(n7257), .A2(prog_data[11]), .B1(\mem[112][11] ), .B2(
        n7256), .Z(n2872) );
  OA22D0 U5017 ( .A1(n7257), .A2(prog_data[10]), .B1(\mem[112][10] ), .B2(
        n7256), .Z(n2871) );
  OA22D0 U5018 ( .A1(n7257), .A2(prog_data[9]), .B1(\mem[112][9] ), .B2(n7256), 
        .Z(n2870) );
  OA22D0 U5019 ( .A1(n7257), .A2(prog_data[8]), .B1(\mem[112][8] ), .B2(n7256), 
        .Z(n2869) );
  OA22D0 U5020 ( .A1(n7257), .A2(prog_data[7]), .B1(\mem[112][7] ), .B2(n7256), 
        .Z(n2868) );
  OA22D0 U5021 ( .A1(n7257), .A2(prog_data[6]), .B1(\mem[112][6] ), .B2(n7256), 
        .Z(n2867) );
  OA22D0 U5022 ( .A1(n7257), .A2(prog_data[5]), .B1(\mem[112][5] ), .B2(n7256), 
        .Z(n2866) );
  OA22D0 U5023 ( .A1(n7257), .A2(prog_data[4]), .B1(\mem[112][4] ), .B2(n7256), 
        .Z(n2865) );
  OA22D0 U5024 ( .A1(n7257), .A2(prog_data[3]), .B1(\mem[112][3] ), .B2(n7256), 
        .Z(n2864) );
  OA22D0 U5025 ( .A1(n7257), .A2(prog_data[2]), .B1(\mem[112][2] ), .B2(n7256), 
        .Z(n2863) );
  OA22D0 U5026 ( .A1(n7257), .A2(prog_data[1]), .B1(\mem[112][1] ), .B2(n7256), 
        .Z(n2862) );
  OA22D0 U5027 ( .A1(n7257), .A2(prog_data[0]), .B1(\mem[112][0] ), .B2(n7256), 
        .Z(n2861) );
  NR2D0 U5028 ( .A1(n7531), .A2(n7286), .ZN(n7258) );
  INVD0 U5029 ( .I(n7258), .ZN(n7259) );
  OA22D0 U5030 ( .A1(n7259), .A2(prog_data[15]), .B1(\mem[113][15] ), .B2(
        n7258), .Z(n2860) );
  OA22D0 U5031 ( .A1(n7259), .A2(prog_data[14]), .B1(\mem[113][14] ), .B2(
        n7258), .Z(n2859) );
  OA22D0 U5032 ( .A1(n7259), .A2(prog_data[13]), .B1(\mem[113][13] ), .B2(
        n7258), .Z(n2858) );
  OA22D0 U5033 ( .A1(n7259), .A2(prog_data[12]), .B1(\mem[113][12] ), .B2(
        n7258), .Z(n2857) );
  OA22D0 U5034 ( .A1(n7259), .A2(prog_data[11]), .B1(\mem[113][11] ), .B2(
        n7258), .Z(n2856) );
  OA22D0 U5035 ( .A1(n7259), .A2(prog_data[10]), .B1(\mem[113][10] ), .B2(
        n7258), .Z(n2855) );
  OA22D0 U5036 ( .A1(n7259), .A2(prog_data[9]), .B1(\mem[113][9] ), .B2(n7258), 
        .Z(n2854) );
  OA22D0 U5037 ( .A1(n7259), .A2(prog_data[8]), .B1(\mem[113][8] ), .B2(n7258), 
        .Z(n2853) );
  OA22D0 U5038 ( .A1(n7259), .A2(prog_data[7]), .B1(\mem[113][7] ), .B2(n7258), 
        .Z(n2852) );
  OA22D0 U5039 ( .A1(n7259), .A2(prog_data[6]), .B1(\mem[113][6] ), .B2(n7258), 
        .Z(n2851) );
  OA22D0 U5040 ( .A1(n7259), .A2(prog_data[5]), .B1(\mem[113][5] ), .B2(n7258), 
        .Z(n2850) );
  OA22D0 U5041 ( .A1(n7259), .A2(prog_data[4]), .B1(\mem[113][4] ), .B2(n7258), 
        .Z(n2849) );
  OA22D0 U5042 ( .A1(n7259), .A2(prog_data[3]), .B1(\mem[113][3] ), .B2(n7258), 
        .Z(n2848) );
  OA22D0 U5043 ( .A1(n7259), .A2(prog_data[2]), .B1(\mem[113][2] ), .B2(n7258), 
        .Z(n2847) );
  OA22D0 U5044 ( .A1(n7259), .A2(prog_data[1]), .B1(\mem[113][1] ), .B2(n7258), 
        .Z(n2846) );
  OA22D0 U5045 ( .A1(n7259), .A2(prog_data[0]), .B1(\mem[113][0] ), .B2(n7258), 
        .Z(n2845) );
  NR2D0 U5046 ( .A1(n7534), .A2(n7286), .ZN(n7260) );
  OA22D0 U5047 ( .A1(n7261), .A2(prog_data[15]), .B1(\mem[114][15] ), .B2(
        n7260), .Z(n2844) );
  OA22D0 U5048 ( .A1(n7261), .A2(prog_data[14]), .B1(\mem[114][14] ), .B2(
        n7260), .Z(n2843) );
  OA22D0 U5049 ( .A1(n7261), .A2(prog_data[13]), .B1(\mem[114][13] ), .B2(
        n7260), .Z(n2842) );
  OA22D0 U5050 ( .A1(n7261), .A2(prog_data[12]), .B1(\mem[114][12] ), .B2(
        n7260), .Z(n2841) );
  OA22D0 U5051 ( .A1(n7261), .A2(prog_data[11]), .B1(\mem[114][11] ), .B2(
        n7260), .Z(n2840) );
  OA22D0 U5052 ( .A1(n7261), .A2(prog_data[10]), .B1(\mem[114][10] ), .B2(
        n7260), .Z(n2839) );
  OA22D0 U5053 ( .A1(n7261), .A2(prog_data[9]), .B1(\mem[114][9] ), .B2(n7260), 
        .Z(n2838) );
  OA22D0 U5054 ( .A1(n7261), .A2(prog_data[8]), .B1(\mem[114][8] ), .B2(n7260), 
        .Z(n2837) );
  OA22D0 U5055 ( .A1(n7261), .A2(prog_data[7]), .B1(\mem[114][7] ), .B2(n7260), 
        .Z(n2836) );
  OA22D0 U5056 ( .A1(n7261), .A2(prog_data[6]), .B1(\mem[114][6] ), .B2(n7260), 
        .Z(n2835) );
  OA22D0 U5057 ( .A1(n7261), .A2(prog_data[5]), .B1(\mem[114][5] ), .B2(n7260), 
        .Z(n2834) );
  OA22D0 U5058 ( .A1(n7261), .A2(prog_data[4]), .B1(\mem[114][4] ), .B2(n7260), 
        .Z(n2833) );
  OA22D0 U5059 ( .A1(n7261), .A2(prog_data[3]), .B1(\mem[114][3] ), .B2(n7260), 
        .Z(n2832) );
  OA22D0 U5060 ( .A1(n7261), .A2(prog_data[2]), .B1(\mem[114][2] ), .B2(n7260), 
        .Z(n2831) );
  OA22D0 U5061 ( .A1(n7261), .A2(prog_data[1]), .B1(\mem[114][1] ), .B2(n7260), 
        .Z(n2830) );
  OA22D0 U5062 ( .A1(n7261), .A2(prog_data[0]), .B1(\mem[114][0] ), .B2(n7260), 
        .Z(n2829) );
  NR2D0 U5063 ( .A1(n7537), .A2(n7286), .ZN(n7262) );
  INVD0 U5064 ( .I(n7262), .ZN(n7263) );
  OA22D0 U5065 ( .A1(n7263), .A2(prog_data[15]), .B1(\mem[115][15] ), .B2(
        n7262), .Z(n2828) );
  OA22D0 U5066 ( .A1(n7263), .A2(prog_data[14]), .B1(\mem[115][14] ), .B2(
        n7262), .Z(n2827) );
  OA22D0 U5067 ( .A1(n7263), .A2(prog_data[13]), .B1(\mem[115][13] ), .B2(
        n7262), .Z(n2826) );
  OA22D0 U5068 ( .A1(n7263), .A2(prog_data[12]), .B1(\mem[115][12] ), .B2(
        n7262), .Z(n2825) );
  OA22D0 U5069 ( .A1(n7263), .A2(prog_data[11]), .B1(\mem[115][11] ), .B2(
        n7262), .Z(n2824) );
  OA22D0 U5070 ( .A1(n7263), .A2(prog_data[10]), .B1(\mem[115][10] ), .B2(
        n7262), .Z(n2823) );
  OA22D0 U5071 ( .A1(n7263), .A2(prog_data[9]), .B1(\mem[115][9] ), .B2(n7262), 
        .Z(n2822) );
  OA22D0 U5072 ( .A1(n7263), .A2(prog_data[8]), .B1(\mem[115][8] ), .B2(n7262), 
        .Z(n2821) );
  OA22D0 U5073 ( .A1(n7263), .A2(prog_data[7]), .B1(\mem[115][7] ), .B2(n7262), 
        .Z(n2820) );
  OA22D0 U5074 ( .A1(n7263), .A2(prog_data[6]), .B1(\mem[115][6] ), .B2(n7262), 
        .Z(n2819) );
  OA22D0 U5075 ( .A1(n7263), .A2(prog_data[5]), .B1(\mem[115][5] ), .B2(n7262), 
        .Z(n2818) );
  OA22D0 U5076 ( .A1(n7263), .A2(prog_data[4]), .B1(\mem[115][4] ), .B2(n7262), 
        .Z(n2817) );
  OA22D0 U5077 ( .A1(n7263), .A2(prog_data[3]), .B1(\mem[115][3] ), .B2(n7262), 
        .Z(n2816) );
  OA22D0 U5078 ( .A1(n7263), .A2(prog_data[2]), .B1(\mem[115][2] ), .B2(n7262), 
        .Z(n2815) );
  OA22D0 U5079 ( .A1(n7263), .A2(prog_data[1]), .B1(\mem[115][1] ), .B2(n7262), 
        .Z(n2814) );
  OA22D0 U5080 ( .A1(n7263), .A2(prog_data[0]), .B1(\mem[115][0] ), .B2(n7262), 
        .Z(n2813) );
  NR2D0 U5081 ( .A1(n7540), .A2(n7286), .ZN(n7264) );
  INVD0 U5082 ( .I(n7264), .ZN(n7265) );
  OA22D0 U5083 ( .A1(n7265), .A2(prog_data[15]), .B1(\mem[116][15] ), .B2(
        n7264), .Z(n2812) );
  OA22D0 U5084 ( .A1(n7265), .A2(prog_data[14]), .B1(\mem[116][14] ), .B2(
        n7264), .Z(n2811) );
  OA22D0 U5085 ( .A1(n7265), .A2(prog_data[13]), .B1(\mem[116][13] ), .B2(
        n7264), .Z(n2810) );
  OA22D0 U5086 ( .A1(n7265), .A2(prog_data[12]), .B1(\mem[116][12] ), .B2(
        n7264), .Z(n2809) );
  OA22D0 U5087 ( .A1(n7265), .A2(prog_data[11]), .B1(\mem[116][11] ), .B2(
        n7264), .Z(n2808) );
  OA22D0 U5088 ( .A1(n7265), .A2(prog_data[10]), .B1(\mem[116][10] ), .B2(
        n7264), .Z(n2807) );
  OA22D0 U5089 ( .A1(n7265), .A2(prog_data[9]), .B1(\mem[116][9] ), .B2(n7264), 
        .Z(n2806) );
  OA22D0 U5090 ( .A1(n7265), .A2(prog_data[8]), .B1(\mem[116][8] ), .B2(n7264), 
        .Z(n2805) );
  OA22D0 U5091 ( .A1(n7265), .A2(prog_data[7]), .B1(\mem[116][7] ), .B2(n7264), 
        .Z(n2804) );
  OA22D0 U5092 ( .A1(n7265), .A2(prog_data[6]), .B1(\mem[116][6] ), .B2(n7264), 
        .Z(n2803) );
  OA22D0 U5093 ( .A1(n7265), .A2(prog_data[5]), .B1(\mem[116][5] ), .B2(n7264), 
        .Z(n2802) );
  OA22D0 U5094 ( .A1(n7265), .A2(prog_data[4]), .B1(\mem[116][4] ), .B2(n7264), 
        .Z(n2801) );
  OA22D0 U5095 ( .A1(n7265), .A2(prog_data[3]), .B1(\mem[116][3] ), .B2(n7264), 
        .Z(n2800) );
  OA22D0 U5096 ( .A1(n7265), .A2(prog_data[2]), .B1(\mem[116][2] ), .B2(n7264), 
        .Z(n2799) );
  OA22D0 U5097 ( .A1(n7265), .A2(prog_data[1]), .B1(\mem[116][1] ), .B2(n7264), 
        .Z(n2798) );
  OA22D0 U5098 ( .A1(n7265), .A2(prog_data[0]), .B1(\mem[116][0] ), .B2(n7264), 
        .Z(n2797) );
  NR2D0 U5099 ( .A1(n7543), .A2(n7286), .ZN(n7266) );
  INVD0 U5100 ( .I(n7266), .ZN(n7267) );
  OA22D0 U5101 ( .A1(n7267), .A2(prog_data[15]), .B1(\mem[117][15] ), .B2(
        n7266), .Z(n2796) );
  OA22D0 U5102 ( .A1(n7267), .A2(prog_data[14]), .B1(\mem[117][14] ), .B2(
        n7266), .Z(n2795) );
  OA22D0 U5103 ( .A1(n7267), .A2(prog_data[13]), .B1(\mem[117][13] ), .B2(
        n7266), .Z(n2794) );
  OA22D0 U5104 ( .A1(n7267), .A2(prog_data[12]), .B1(\mem[117][12] ), .B2(
        n7266), .Z(n2793) );
  OA22D0 U5105 ( .A1(n7267), .A2(prog_data[11]), .B1(\mem[117][11] ), .B2(
        n7266), .Z(n2792) );
  OA22D0 U5106 ( .A1(n7267), .A2(prog_data[10]), .B1(\mem[117][10] ), .B2(
        n7266), .Z(n2791) );
  OA22D0 U5107 ( .A1(n7267), .A2(prog_data[9]), .B1(\mem[117][9] ), .B2(n7266), 
        .Z(n2790) );
  OA22D0 U5108 ( .A1(n7267), .A2(prog_data[8]), .B1(\mem[117][8] ), .B2(n7266), 
        .Z(n2789) );
  OA22D0 U5109 ( .A1(n7267), .A2(prog_data[7]), .B1(\mem[117][7] ), .B2(n7266), 
        .Z(n2788) );
  OA22D0 U5110 ( .A1(n7267), .A2(prog_data[6]), .B1(\mem[117][6] ), .B2(n7266), 
        .Z(n2787) );
  OA22D0 U5111 ( .A1(n7267), .A2(prog_data[5]), .B1(\mem[117][5] ), .B2(n7266), 
        .Z(n2786) );
  OA22D0 U5112 ( .A1(n7267), .A2(prog_data[4]), .B1(\mem[117][4] ), .B2(n7266), 
        .Z(n2785) );
  OA22D0 U5113 ( .A1(n7267), .A2(prog_data[3]), .B1(\mem[117][3] ), .B2(n7266), 
        .Z(n2784) );
  OA22D0 U5114 ( .A1(n7267), .A2(prog_data[2]), .B1(\mem[117][2] ), .B2(n7266), 
        .Z(n2783) );
  OA22D0 U5115 ( .A1(n7267), .A2(prog_data[1]), .B1(\mem[117][1] ), .B2(n7266), 
        .Z(n2782) );
  OA22D0 U5116 ( .A1(n7267), .A2(prog_data[0]), .B1(\mem[117][0] ), .B2(n7266), 
        .Z(n2781) );
  NR2D0 U5117 ( .A1(n7546), .A2(n7286), .ZN(n7268) );
  INVD0 U5118 ( .I(n7268), .ZN(n7269) );
  OA22D0 U5119 ( .A1(n7269), .A2(prog_data[15]), .B1(\mem[118][15] ), .B2(
        n7268), .Z(n2780) );
  OA22D0 U5120 ( .A1(n7269), .A2(prog_data[14]), .B1(\mem[118][14] ), .B2(
        n7268), .Z(n2779) );
  OA22D0 U5121 ( .A1(n7269), .A2(prog_data[13]), .B1(\mem[118][13] ), .B2(
        n7268), .Z(n2778) );
  OA22D0 U5122 ( .A1(n7269), .A2(prog_data[12]), .B1(\mem[118][12] ), .B2(
        n7268), .Z(n2777) );
  OA22D0 U5123 ( .A1(n7269), .A2(prog_data[11]), .B1(\mem[118][11] ), .B2(
        n7268), .Z(n2776) );
  OA22D0 U5124 ( .A1(n7269), .A2(prog_data[10]), .B1(\mem[118][10] ), .B2(
        n7268), .Z(n2775) );
  OA22D0 U5125 ( .A1(n7269), .A2(prog_data[9]), .B1(\mem[118][9] ), .B2(n7268), 
        .Z(n2774) );
  OA22D0 U5126 ( .A1(n7269), .A2(prog_data[8]), .B1(\mem[118][8] ), .B2(n7268), 
        .Z(n2773) );
  OA22D0 U5127 ( .A1(n7269), .A2(prog_data[7]), .B1(\mem[118][7] ), .B2(n7268), 
        .Z(n2772) );
  OA22D0 U5128 ( .A1(n7269), .A2(prog_data[6]), .B1(\mem[118][6] ), .B2(n7268), 
        .Z(n2771) );
  OA22D0 U5129 ( .A1(n7269), .A2(prog_data[5]), .B1(\mem[118][5] ), .B2(n7268), 
        .Z(n2770) );
  OA22D0 U5130 ( .A1(n7269), .A2(prog_data[4]), .B1(\mem[118][4] ), .B2(n7268), 
        .Z(n2769) );
  OA22D0 U5131 ( .A1(n7269), .A2(prog_data[3]), .B1(\mem[118][3] ), .B2(n7268), 
        .Z(n2768) );
  OA22D0 U5132 ( .A1(n7269), .A2(prog_data[2]), .B1(\mem[118][2] ), .B2(n7268), 
        .Z(n2767) );
  OA22D0 U5133 ( .A1(n7269), .A2(prog_data[1]), .B1(\mem[118][1] ), .B2(n7268), 
        .Z(n2766) );
  OA22D0 U5134 ( .A1(n7269), .A2(prog_data[0]), .B1(\mem[118][0] ), .B2(n7268), 
        .Z(n2765) );
  NR2D0 U5135 ( .A1(n7549), .A2(n7286), .ZN(n7270) );
  INVD0 U5136 ( .I(n7270), .ZN(n7271) );
  OA22D0 U5137 ( .A1(n7271), .A2(prog_data[15]), .B1(\mem[119][15] ), .B2(
        n7270), .Z(n2764) );
  OA22D0 U5138 ( .A1(n7271), .A2(prog_data[14]), .B1(\mem[119][14] ), .B2(
        n7270), .Z(n2763) );
  OA22D0 U5139 ( .A1(n7271), .A2(prog_data[13]), .B1(\mem[119][13] ), .B2(
        n7270), .Z(n2762) );
  OA22D0 U5140 ( .A1(n7271), .A2(prog_data[12]), .B1(\mem[119][12] ), .B2(
        n7270), .Z(n2761) );
  OA22D0 U5141 ( .A1(n7271), .A2(prog_data[11]), .B1(\mem[119][11] ), .B2(
        n7270), .Z(n2760) );
  OA22D0 U5142 ( .A1(n7271), .A2(prog_data[10]), .B1(\mem[119][10] ), .B2(
        n7270), .Z(n2759) );
  OA22D0 U5143 ( .A1(n7271), .A2(prog_data[9]), .B1(\mem[119][9] ), .B2(n7270), 
        .Z(n2758) );
  OA22D0 U5144 ( .A1(n7271), .A2(prog_data[8]), .B1(\mem[119][8] ), .B2(n7270), 
        .Z(n2757) );
  OA22D0 U5145 ( .A1(n7271), .A2(prog_data[7]), .B1(\mem[119][7] ), .B2(n7270), 
        .Z(n2756) );
  OA22D0 U5146 ( .A1(n7271), .A2(prog_data[6]), .B1(\mem[119][6] ), .B2(n7270), 
        .Z(n2755) );
  OA22D0 U5147 ( .A1(n7271), .A2(prog_data[5]), .B1(\mem[119][5] ), .B2(n7270), 
        .Z(n2754) );
  OA22D0 U5148 ( .A1(n7271), .A2(prog_data[4]), .B1(\mem[119][4] ), .B2(n7270), 
        .Z(n2753) );
  OA22D0 U5149 ( .A1(n7271), .A2(prog_data[3]), .B1(\mem[119][3] ), .B2(n7270), 
        .Z(n2752) );
  OA22D0 U5150 ( .A1(n7271), .A2(prog_data[2]), .B1(\mem[119][2] ), .B2(n7270), 
        .Z(n2751) );
  OA22D0 U5151 ( .A1(n7271), .A2(prog_data[1]), .B1(\mem[119][1] ), .B2(n7270), 
        .Z(n2750) );
  OA22D0 U5152 ( .A1(n7271), .A2(prog_data[0]), .B1(\mem[119][0] ), .B2(n7270), 
        .Z(n2749) );
  NR2D0 U5153 ( .A1(n7552), .A2(n7286), .ZN(n7272) );
  INVD0 U5154 ( .I(n7272), .ZN(n7273) );
  OA22D0 U5155 ( .A1(n7273), .A2(prog_data[15]), .B1(\mem[120][15] ), .B2(
        n7272), .Z(n2748) );
  OA22D0 U5156 ( .A1(n7273), .A2(prog_data[14]), .B1(\mem[120][14] ), .B2(
        n7272), .Z(n2747) );
  OA22D0 U5157 ( .A1(n7273), .A2(prog_data[13]), .B1(\mem[120][13] ), .B2(
        n7272), .Z(n2746) );
  OA22D0 U5158 ( .A1(n7273), .A2(prog_data[12]), .B1(\mem[120][12] ), .B2(
        n7272), .Z(n2745) );
  OA22D0 U5159 ( .A1(n7273), .A2(prog_data[11]), .B1(\mem[120][11] ), .B2(
        n7272), .Z(n2744) );
  OA22D0 U5160 ( .A1(n7273), .A2(prog_data[10]), .B1(\mem[120][10] ), .B2(
        n7272), .Z(n2743) );
  OA22D0 U5161 ( .A1(n7273), .A2(prog_data[9]), .B1(\mem[120][9] ), .B2(n7272), 
        .Z(n2742) );
  OA22D0 U5162 ( .A1(n7273), .A2(prog_data[8]), .B1(\mem[120][8] ), .B2(n7272), 
        .Z(n2741) );
  OA22D0 U5163 ( .A1(n7273), .A2(prog_data[7]), .B1(\mem[120][7] ), .B2(n7272), 
        .Z(n2740) );
  OA22D0 U5164 ( .A1(n7273), .A2(prog_data[6]), .B1(\mem[120][6] ), .B2(n7272), 
        .Z(n2739) );
  OA22D0 U5165 ( .A1(n7273), .A2(prog_data[5]), .B1(\mem[120][5] ), .B2(n7272), 
        .Z(n2738) );
  OA22D0 U5166 ( .A1(n7273), .A2(prog_data[4]), .B1(\mem[120][4] ), .B2(n7272), 
        .Z(n2737) );
  OA22D0 U5167 ( .A1(n7273), .A2(prog_data[3]), .B1(\mem[120][3] ), .B2(n7272), 
        .Z(n2736) );
  OA22D0 U5168 ( .A1(n7273), .A2(prog_data[2]), .B1(\mem[120][2] ), .B2(n7272), 
        .Z(n2735) );
  OA22D0 U5169 ( .A1(n7273), .A2(prog_data[1]), .B1(\mem[120][1] ), .B2(n7272), 
        .Z(n2734) );
  OA22D0 U5170 ( .A1(n7273), .A2(prog_data[0]), .B1(\mem[120][0] ), .B2(n7272), 
        .Z(n2733) );
  INVD0 U5171 ( .I(n7274), .ZN(n7275) );
  OA22D0 U5172 ( .A1(n7275), .A2(prog_data[15]), .B1(\mem[121][15] ), .B2(
        n7274), .Z(n2732) );
  OA22D0 U5173 ( .A1(n7275), .A2(prog_data[14]), .B1(\mem[121][14] ), .B2(
        n7274), .Z(n2731) );
  OA22D0 U5174 ( .A1(n7275), .A2(prog_data[13]), .B1(\mem[121][13] ), .B2(
        n7274), .Z(n2730) );
  OA22D0 U5175 ( .A1(n7275), .A2(prog_data[12]), .B1(\mem[121][12] ), .B2(
        n7274), .Z(n2729) );
  OA22D0 U5176 ( .A1(n7275), .A2(prog_data[11]), .B1(\mem[121][11] ), .B2(
        n7274), .Z(n2728) );
  OA22D0 U5177 ( .A1(n7275), .A2(prog_data[10]), .B1(\mem[121][10] ), .B2(
        n7274), .Z(n2727) );
  OA22D0 U5178 ( .A1(n7275), .A2(prog_data[9]), .B1(\mem[121][9] ), .B2(n7274), 
        .Z(n2726) );
  OA22D0 U5179 ( .A1(n7275), .A2(prog_data[8]), .B1(\mem[121][8] ), .B2(n7274), 
        .Z(n2725) );
  OA22D0 U5180 ( .A1(n7275), .A2(prog_data[7]), .B1(\mem[121][7] ), .B2(n7274), 
        .Z(n2724) );
  OA22D0 U5181 ( .A1(n7275), .A2(prog_data[6]), .B1(\mem[121][6] ), .B2(n7274), 
        .Z(n2723) );
  OA22D0 U5182 ( .A1(n7275), .A2(prog_data[5]), .B1(\mem[121][5] ), .B2(n7274), 
        .Z(n2722) );
  OA22D0 U5183 ( .A1(n7275), .A2(prog_data[4]), .B1(\mem[121][4] ), .B2(n7274), 
        .Z(n2721) );
  OA22D0 U5184 ( .A1(n7275), .A2(prog_data[3]), .B1(\mem[121][3] ), .B2(n7274), 
        .Z(n2720) );
  OA22D0 U5185 ( .A1(n7275), .A2(prog_data[2]), .B1(\mem[121][2] ), .B2(n7274), 
        .Z(n2719) );
  OA22D0 U5186 ( .A1(n7275), .A2(prog_data[1]), .B1(\mem[121][1] ), .B2(n7274), 
        .Z(n2718) );
  OA22D0 U5187 ( .A1(n7275), .A2(prog_data[0]), .B1(\mem[121][0] ), .B2(n7274), 
        .Z(n2717) );
  NR2D0 U5188 ( .A1(n7558), .A2(n7286), .ZN(n7276) );
  INVD0 U5189 ( .I(n7276), .ZN(n7277) );
  OA22D0 U5190 ( .A1(n7277), .A2(prog_data[15]), .B1(\mem[122][15] ), .B2(
        n7276), .Z(n2716) );
  OA22D0 U5191 ( .A1(n7277), .A2(prog_data[14]), .B1(\mem[122][14] ), .B2(
        n7276), .Z(n2715) );
  OA22D0 U5192 ( .A1(n7277), .A2(prog_data[13]), .B1(\mem[122][13] ), .B2(
        n7276), .Z(n2714) );
  OA22D0 U5193 ( .A1(n7277), .A2(prog_data[12]), .B1(\mem[122][12] ), .B2(
        n7276), .Z(n2713) );
  OA22D0 U5194 ( .A1(n7277), .A2(prog_data[11]), .B1(\mem[122][11] ), .B2(
        n7276), .Z(n2712) );
  OA22D0 U5195 ( .A1(n7277), .A2(prog_data[10]), .B1(\mem[122][10] ), .B2(
        n7276), .Z(n2711) );
  OA22D0 U5196 ( .A1(n7277), .A2(prog_data[9]), .B1(\mem[122][9] ), .B2(n7276), 
        .Z(n2710) );
  OA22D0 U5197 ( .A1(n7277), .A2(prog_data[8]), .B1(\mem[122][8] ), .B2(n7276), 
        .Z(n2709) );
  OA22D0 U5198 ( .A1(n7277), .A2(prog_data[7]), .B1(\mem[122][7] ), .B2(n7276), 
        .Z(n2708) );
  OA22D0 U5199 ( .A1(n7277), .A2(prog_data[6]), .B1(\mem[122][6] ), .B2(n7276), 
        .Z(n2707) );
  OA22D0 U5200 ( .A1(n7277), .A2(prog_data[5]), .B1(\mem[122][5] ), .B2(n7276), 
        .Z(n2706) );
  OA22D0 U5201 ( .A1(n7277), .A2(prog_data[4]), .B1(\mem[122][4] ), .B2(n7276), 
        .Z(n2705) );
  OA22D0 U5202 ( .A1(n7277), .A2(prog_data[3]), .B1(\mem[122][3] ), .B2(n7276), 
        .Z(n2704) );
  OA22D0 U5203 ( .A1(n7277), .A2(prog_data[2]), .B1(\mem[122][2] ), .B2(n7276), 
        .Z(n2703) );
  OA22D0 U5204 ( .A1(n7277), .A2(prog_data[1]), .B1(\mem[122][1] ), .B2(n7276), 
        .Z(n2702) );
  OA22D0 U5205 ( .A1(n7277), .A2(prog_data[0]), .B1(\mem[122][0] ), .B2(n7276), 
        .Z(n2701) );
  NR2D0 U5206 ( .A1(n7561), .A2(n7286), .ZN(n7278) );
  INVD0 U5207 ( .I(n7278), .ZN(n7279) );
  OA22D0 U5208 ( .A1(n7279), .A2(prog_data[15]), .B1(\mem[123][15] ), .B2(
        n7278), .Z(n2700) );
  OA22D0 U5209 ( .A1(n7279), .A2(prog_data[14]), .B1(\mem[123][14] ), .B2(
        n7278), .Z(n2699) );
  OA22D0 U5210 ( .A1(n7279), .A2(prog_data[13]), .B1(\mem[123][13] ), .B2(
        n7278), .Z(n2698) );
  OA22D0 U5211 ( .A1(n7279), .A2(prog_data[12]), .B1(\mem[123][12] ), .B2(
        n7278), .Z(n2697) );
  OA22D0 U5212 ( .A1(n7279), .A2(prog_data[11]), .B1(\mem[123][11] ), .B2(
        n7278), .Z(n2696) );
  OA22D0 U5213 ( .A1(n7279), .A2(prog_data[10]), .B1(\mem[123][10] ), .B2(
        n7278), .Z(n2695) );
  OA22D0 U5214 ( .A1(n7279), .A2(prog_data[9]), .B1(\mem[123][9] ), .B2(n7278), 
        .Z(n2694) );
  OA22D0 U5215 ( .A1(n7279), .A2(prog_data[8]), .B1(\mem[123][8] ), .B2(n7278), 
        .Z(n2693) );
  OA22D0 U5216 ( .A1(n7279), .A2(prog_data[7]), .B1(\mem[123][7] ), .B2(n7278), 
        .Z(n2692) );
  OA22D0 U5217 ( .A1(n7279), .A2(prog_data[6]), .B1(\mem[123][6] ), .B2(n7278), 
        .Z(n2691) );
  OA22D0 U5218 ( .A1(n7279), .A2(prog_data[5]), .B1(\mem[123][5] ), .B2(n7278), 
        .Z(n2690) );
  OA22D0 U5219 ( .A1(n7279), .A2(prog_data[4]), .B1(\mem[123][4] ), .B2(n7278), 
        .Z(n2689) );
  OA22D0 U5220 ( .A1(n7279), .A2(prog_data[3]), .B1(\mem[123][3] ), .B2(n7278), 
        .Z(n2688) );
  OA22D0 U5221 ( .A1(n7279), .A2(prog_data[2]), .B1(\mem[123][2] ), .B2(n7278), 
        .Z(n2687) );
  OA22D0 U5222 ( .A1(n7279), .A2(prog_data[1]), .B1(\mem[123][1] ), .B2(n7278), 
        .Z(n2686) );
  OA22D0 U5223 ( .A1(n7279), .A2(prog_data[0]), .B1(\mem[123][0] ), .B2(n7278), 
        .Z(n2685) );
  NR2D0 U5224 ( .A1(n7564), .A2(n7286), .ZN(n7280) );
  INVD0 U5225 ( .I(n7280), .ZN(n7281) );
  OA22D0 U5226 ( .A1(n7281), .A2(prog_data[15]), .B1(\mem[124][15] ), .B2(
        n7280), .Z(n2684) );
  OA22D0 U5227 ( .A1(n7281), .A2(prog_data[14]), .B1(\mem[124][14] ), .B2(
        n7280), .Z(n2683) );
  OA22D0 U5228 ( .A1(n7281), .A2(prog_data[13]), .B1(\mem[124][13] ), .B2(
        n7280), .Z(n2682) );
  OA22D0 U5229 ( .A1(n7281), .A2(prog_data[12]), .B1(\mem[124][12] ), .B2(
        n7280), .Z(n2681) );
  OA22D0 U5230 ( .A1(n7281), .A2(prog_data[11]), .B1(\mem[124][11] ), .B2(
        n7280), .Z(n2680) );
  OA22D0 U5231 ( .A1(n7281), .A2(prog_data[10]), .B1(\mem[124][10] ), .B2(
        n7280), .Z(n2679) );
  OA22D0 U5232 ( .A1(n7281), .A2(prog_data[9]), .B1(\mem[124][9] ), .B2(n7280), 
        .Z(n2678) );
  OA22D0 U5233 ( .A1(n7281), .A2(prog_data[8]), .B1(\mem[124][8] ), .B2(n7280), 
        .Z(n2677) );
  OA22D0 U5234 ( .A1(n7281), .A2(prog_data[7]), .B1(\mem[124][7] ), .B2(n7280), 
        .Z(n2676) );
  OA22D0 U5235 ( .A1(n7281), .A2(prog_data[6]), .B1(\mem[124][6] ), .B2(n7280), 
        .Z(n2675) );
  OA22D0 U5236 ( .A1(n7281), .A2(prog_data[5]), .B1(\mem[124][5] ), .B2(n7280), 
        .Z(n2674) );
  OA22D0 U5237 ( .A1(n7281), .A2(prog_data[4]), .B1(\mem[124][4] ), .B2(n7280), 
        .Z(n2673) );
  OA22D0 U5238 ( .A1(n7281), .A2(prog_data[3]), .B1(\mem[124][3] ), .B2(n7280), 
        .Z(n2672) );
  OA22D0 U5239 ( .A1(n7281), .A2(prog_data[2]), .B1(\mem[124][2] ), .B2(n7280), 
        .Z(n2671) );
  OA22D0 U5240 ( .A1(n7281), .A2(prog_data[1]), .B1(\mem[124][1] ), .B2(n7280), 
        .Z(n2670) );
  OA22D0 U5241 ( .A1(n7281), .A2(prog_data[0]), .B1(\mem[124][0] ), .B2(n7280), 
        .Z(n2669) );
  NR2D0 U5242 ( .A1(n7567), .A2(n7286), .ZN(n7282) );
  INVD0 U5243 ( .I(n7282), .ZN(n7283) );
  OA22D0 U5244 ( .A1(n7283), .A2(prog_data[15]), .B1(\mem[125][15] ), .B2(
        n7282), .Z(n2668) );
  OA22D0 U5245 ( .A1(n7283), .A2(prog_data[14]), .B1(\mem[125][14] ), .B2(
        n7282), .Z(n2667) );
  OA22D0 U5246 ( .A1(n7283), .A2(prog_data[13]), .B1(\mem[125][13] ), .B2(
        n7282), .Z(n2666) );
  OA22D0 U5247 ( .A1(n7283), .A2(prog_data[12]), .B1(\mem[125][12] ), .B2(
        n7282), .Z(n2665) );
  OA22D0 U5248 ( .A1(n7283), .A2(prog_data[11]), .B1(\mem[125][11] ), .B2(
        n7282), .Z(n2664) );
  OA22D0 U5249 ( .A1(n7283), .A2(prog_data[10]), .B1(\mem[125][10] ), .B2(
        n7282), .Z(n2663) );
  OA22D0 U5250 ( .A1(n7283), .A2(prog_data[9]), .B1(\mem[125][9] ), .B2(n7282), 
        .Z(n2662) );
  OA22D0 U5251 ( .A1(n7283), .A2(prog_data[8]), .B1(\mem[125][8] ), .B2(n7282), 
        .Z(n2661) );
  OA22D0 U5252 ( .A1(n7283), .A2(prog_data[7]), .B1(\mem[125][7] ), .B2(n7282), 
        .Z(n2660) );
  OA22D0 U5253 ( .A1(n7283), .A2(prog_data[6]), .B1(\mem[125][6] ), .B2(n7282), 
        .Z(n2659) );
  OA22D0 U5254 ( .A1(n7283), .A2(prog_data[5]), .B1(\mem[125][5] ), .B2(n7282), 
        .Z(n2658) );
  OA22D0 U5255 ( .A1(n7283), .A2(prog_data[4]), .B1(\mem[125][4] ), .B2(n7282), 
        .Z(n2657) );
  OA22D0 U5256 ( .A1(n7283), .A2(prog_data[3]), .B1(\mem[125][3] ), .B2(n7282), 
        .Z(n2656) );
  OA22D0 U5257 ( .A1(n7283), .A2(prog_data[2]), .B1(\mem[125][2] ), .B2(n7282), 
        .Z(n2655) );
  OA22D0 U5258 ( .A1(n7283), .A2(prog_data[1]), .B1(\mem[125][1] ), .B2(n7282), 
        .Z(n2654) );
  OA22D0 U5259 ( .A1(n7283), .A2(prog_data[0]), .B1(\mem[125][0] ), .B2(n7282), 
        .Z(n2653) );
  NR2D0 U5260 ( .A1(n7570), .A2(n7286), .ZN(n7284) );
  INVD0 U5261 ( .I(n7284), .ZN(n7285) );
  OA22D0 U5262 ( .A1(n7285), .A2(prog_data[15]), .B1(\mem[126][15] ), .B2(
        n7284), .Z(n2652) );
  OA22D0 U5263 ( .A1(n7285), .A2(prog_data[14]), .B1(\mem[126][14] ), .B2(
        n7284), .Z(n2651) );
  OA22D0 U5264 ( .A1(n7285), .A2(prog_data[13]), .B1(\mem[126][13] ), .B2(
        n7284), .Z(n2650) );
  OA22D0 U5265 ( .A1(n7285), .A2(prog_data[12]), .B1(\mem[126][12] ), .B2(
        n7284), .Z(n2649) );
  OA22D0 U5266 ( .A1(n7285), .A2(prog_data[11]), .B1(\mem[126][11] ), .B2(
        n7284), .Z(n2648) );
  OA22D0 U5267 ( .A1(n7285), .A2(prog_data[10]), .B1(\mem[126][10] ), .B2(
        n7284), .Z(n2647) );
  OA22D0 U5268 ( .A1(n7285), .A2(prog_data[9]), .B1(\mem[126][9] ), .B2(n7284), 
        .Z(n2646) );
  OA22D0 U5269 ( .A1(n7285), .A2(prog_data[8]), .B1(\mem[126][8] ), .B2(n7284), 
        .Z(n2645) );
  OA22D0 U5270 ( .A1(n7285), .A2(prog_data[7]), .B1(\mem[126][7] ), .B2(n7284), 
        .Z(n2644) );
  OA22D0 U5271 ( .A1(n7285), .A2(prog_data[6]), .B1(\mem[126][6] ), .B2(n7284), 
        .Z(n2643) );
  OA22D0 U5272 ( .A1(n7285), .A2(prog_data[5]), .B1(\mem[126][5] ), .B2(n7284), 
        .Z(n2642) );
  OA22D0 U5273 ( .A1(n7285), .A2(prog_data[4]), .B1(\mem[126][4] ), .B2(n7284), 
        .Z(n2641) );
  OA22D0 U5274 ( .A1(n7285), .A2(prog_data[3]), .B1(\mem[126][3] ), .B2(n7284), 
        .Z(n2640) );
  OA22D0 U5275 ( .A1(n7285), .A2(prog_data[2]), .B1(\mem[126][2] ), .B2(n7284), 
        .Z(n2639) );
  OA22D0 U5276 ( .A1(n7285), .A2(prog_data[1]), .B1(\mem[126][1] ), .B2(n7284), 
        .Z(n2638) );
  OA22D0 U5277 ( .A1(n7285), .A2(prog_data[0]), .B1(\mem[126][0] ), .B2(n7284), 
        .Z(n2637) );
  NR2D0 U5278 ( .A1(n7574), .A2(n7286), .ZN(n7287) );
  INVD0 U5279 ( .I(n7287), .ZN(n7288) );
  OA22D0 U5280 ( .A1(n7288), .A2(prog_data[15]), .B1(\mem[127][15] ), .B2(
        n7287), .Z(n2636) );
  OA22D0 U5281 ( .A1(n7288), .A2(prog_data[14]), .B1(\mem[127][14] ), .B2(
        n7287), .Z(n2635) );
  OA22D0 U5282 ( .A1(n7288), .A2(prog_data[13]), .B1(\mem[127][13] ), .B2(
        n7287), .Z(n2634) );
  OA22D0 U5283 ( .A1(n7288), .A2(prog_data[12]), .B1(\mem[127][12] ), .B2(
        n7287), .Z(n2633) );
  OA22D0 U5284 ( .A1(n7288), .A2(prog_data[11]), .B1(\mem[127][11] ), .B2(
        n7287), .Z(n2632) );
  OA22D0 U5285 ( .A1(n7288), .A2(prog_data[10]), .B1(\mem[127][10] ), .B2(
        n7287), .Z(n2631) );
  OA22D0 U5286 ( .A1(n7288), .A2(prog_data[9]), .B1(\mem[127][9] ), .B2(n7287), 
        .Z(n2630) );
  OA22D0 U5287 ( .A1(n7288), .A2(prog_data[8]), .B1(\mem[127][8] ), .B2(n7287), 
        .Z(n2629) );
  OA22D0 U5288 ( .A1(n7288), .A2(prog_data[7]), .B1(\mem[127][7] ), .B2(n7287), 
        .Z(n2628) );
  OA22D0 U5289 ( .A1(n7288), .A2(prog_data[6]), .B1(\mem[127][6] ), .B2(n7287), 
        .Z(n2627) );
  OA22D0 U5290 ( .A1(n7288), .A2(prog_data[5]), .B1(\mem[127][5] ), .B2(n7287), 
        .Z(n2626) );
  OA22D0 U5291 ( .A1(n7288), .A2(prog_data[4]), .B1(\mem[127][4] ), .B2(n7287), 
        .Z(n2625) );
  OA22D0 U5292 ( .A1(n7288), .A2(prog_data[3]), .B1(\mem[127][3] ), .B2(n7287), 
        .Z(n2624) );
  OA22D0 U5293 ( .A1(n7288), .A2(prog_data[2]), .B1(\mem[127][2] ), .B2(n7287), 
        .Z(n2623) );
  OA22D0 U5294 ( .A1(n7288), .A2(prog_data[1]), .B1(\mem[127][1] ), .B2(n7287), 
        .Z(n2622) );
  OA22D0 U5295 ( .A1(n7288), .A2(prog_data[0]), .B1(\mem[127][0] ), .B2(n7287), 
        .Z(n2621) );
  NR2D0 U5296 ( .A1(prog_addr[4]), .A2(n7322), .ZN(n7492) );
  CKND2D0 U5297 ( .A1(n7324), .A2(n7492), .ZN(n7319) );
  NR2D0 U5298 ( .A1(n7528), .A2(n7319), .ZN(n7289) );
  INVD0 U5299 ( .I(n7289), .ZN(n7290) );
  OA22D0 U5300 ( .A1(n7290), .A2(prog_data[15]), .B1(\mem[128][15] ), .B2(
        n7289), .Z(n2620) );
  OA22D0 U5301 ( .A1(n7290), .A2(prog_data[14]), .B1(\mem[128][14] ), .B2(
        n7289), .Z(n2619) );
  OA22D0 U5302 ( .A1(n7290), .A2(prog_data[13]), .B1(\mem[128][13] ), .B2(
        n7289), .Z(n2618) );
  OA22D0 U5303 ( .A1(n7290), .A2(prog_data[12]), .B1(\mem[128][12] ), .B2(
        n7289), .Z(n2617) );
  OA22D0 U5304 ( .A1(n7290), .A2(prog_data[11]), .B1(\mem[128][11] ), .B2(
        n7289), .Z(n2616) );
  OA22D0 U5305 ( .A1(n7290), .A2(prog_data[10]), .B1(\mem[128][10] ), .B2(
        n7289), .Z(n2615) );
  OA22D0 U5306 ( .A1(n7290), .A2(prog_data[9]), .B1(\mem[128][9] ), .B2(n7289), 
        .Z(n2614) );
  OA22D0 U5307 ( .A1(n7290), .A2(prog_data[8]), .B1(\mem[128][8] ), .B2(n7289), 
        .Z(n2613) );
  OA22D0 U5308 ( .A1(n7290), .A2(prog_data[7]), .B1(\mem[128][7] ), .B2(n7289), 
        .Z(n2612) );
  OA22D0 U5309 ( .A1(n7290), .A2(prog_data[6]), .B1(\mem[128][6] ), .B2(n7289), 
        .Z(n2611) );
  OA22D0 U5310 ( .A1(n7290), .A2(prog_data[5]), .B1(\mem[128][5] ), .B2(n7289), 
        .Z(n2610) );
  OA22D0 U5311 ( .A1(n7290), .A2(prog_data[4]), .B1(\mem[128][4] ), .B2(n7289), 
        .Z(n2609) );
  OA22D0 U5312 ( .A1(n7290), .A2(prog_data[3]), .B1(\mem[128][3] ), .B2(n7289), 
        .Z(n2608) );
  OA22D0 U5313 ( .A1(n7290), .A2(prog_data[2]), .B1(\mem[128][2] ), .B2(n7289), 
        .Z(n2607) );
  OA22D0 U5314 ( .A1(n7290), .A2(prog_data[1]), .B1(\mem[128][1] ), .B2(n7289), 
        .Z(n2606) );
  OA22D0 U5315 ( .A1(n7290), .A2(prog_data[0]), .B1(\mem[128][0] ), .B2(n7289), 
        .Z(n2605) );
  NR2D0 U5316 ( .A1(n7531), .A2(n7319), .ZN(n7291) );
  OA22D0 U5317 ( .A1(n7292), .A2(prog_data[15]), .B1(\mem[129][15] ), .B2(
        n7291), .Z(n2604) );
  OA22D0 U5318 ( .A1(n7292), .A2(prog_data[14]), .B1(\mem[129][14] ), .B2(
        n7291), .Z(n2603) );
  OA22D0 U5319 ( .A1(n7292), .A2(prog_data[13]), .B1(\mem[129][13] ), .B2(
        n7291), .Z(n2602) );
  OA22D0 U5320 ( .A1(n7292), .A2(prog_data[12]), .B1(\mem[129][12] ), .B2(
        n7291), .Z(n2601) );
  OA22D0 U5321 ( .A1(n7292), .A2(prog_data[11]), .B1(\mem[129][11] ), .B2(
        n7291), .Z(n2600) );
  OA22D0 U5322 ( .A1(n7292), .A2(prog_data[10]), .B1(\mem[129][10] ), .B2(
        n7291), .Z(n2599) );
  OA22D0 U5323 ( .A1(n7292), .A2(prog_data[9]), .B1(\mem[129][9] ), .B2(n7291), 
        .Z(n2598) );
  OA22D0 U5324 ( .A1(n7292), .A2(prog_data[8]), .B1(\mem[129][8] ), .B2(n7291), 
        .Z(n2597) );
  OA22D0 U5325 ( .A1(n7292), .A2(prog_data[7]), .B1(\mem[129][7] ), .B2(n7291), 
        .Z(n2596) );
  OA22D0 U5326 ( .A1(n7292), .A2(prog_data[6]), .B1(\mem[129][6] ), .B2(n7291), 
        .Z(n2595) );
  OA22D0 U5327 ( .A1(n7292), .A2(prog_data[5]), .B1(\mem[129][5] ), .B2(n7291), 
        .Z(n2594) );
  OA22D0 U5328 ( .A1(n7292), .A2(prog_data[4]), .B1(\mem[129][4] ), .B2(n7291), 
        .Z(n2593) );
  OA22D0 U5329 ( .A1(n7292), .A2(prog_data[3]), .B1(\mem[129][3] ), .B2(n7291), 
        .Z(n2592) );
  OA22D0 U5330 ( .A1(n7292), .A2(prog_data[2]), .B1(\mem[129][2] ), .B2(n7291), 
        .Z(n2591) );
  OA22D0 U5331 ( .A1(n7292), .A2(prog_data[1]), .B1(\mem[129][1] ), .B2(n7291), 
        .Z(n2590) );
  OA22D0 U5332 ( .A1(n7292), .A2(prog_data[0]), .B1(\mem[129][0] ), .B2(n7291), 
        .Z(n2589) );
  NR2D0 U5333 ( .A1(n7534), .A2(n7319), .ZN(n7293) );
  INVD0 U5334 ( .I(n7293), .ZN(n7294) );
  OA22D0 U5335 ( .A1(n7294), .A2(prog_data[15]), .B1(\mem[130][15] ), .B2(
        n7293), .Z(n2588) );
  OA22D0 U5336 ( .A1(n7294), .A2(prog_data[14]), .B1(\mem[130][14] ), .B2(
        n7293), .Z(n2587) );
  OA22D0 U5337 ( .A1(n7294), .A2(prog_data[13]), .B1(\mem[130][13] ), .B2(
        n7293), .Z(n2586) );
  OA22D0 U5338 ( .A1(n7294), .A2(prog_data[12]), .B1(\mem[130][12] ), .B2(
        n7293), .Z(n2585) );
  OA22D0 U5339 ( .A1(n7294), .A2(prog_data[11]), .B1(\mem[130][11] ), .B2(
        n7293), .Z(n2584) );
  OA22D0 U5340 ( .A1(n7294), .A2(prog_data[10]), .B1(\mem[130][10] ), .B2(
        n7293), .Z(n2583) );
  OA22D0 U5341 ( .A1(n7294), .A2(prog_data[9]), .B1(\mem[130][9] ), .B2(n7293), 
        .Z(n2582) );
  OA22D0 U5342 ( .A1(n7294), .A2(prog_data[8]), .B1(\mem[130][8] ), .B2(n7293), 
        .Z(n2581) );
  OA22D0 U5343 ( .A1(n7294), .A2(prog_data[7]), .B1(\mem[130][7] ), .B2(n7293), 
        .Z(n2580) );
  OA22D0 U5344 ( .A1(n7294), .A2(prog_data[6]), .B1(\mem[130][6] ), .B2(n7293), 
        .Z(n2579) );
  OA22D0 U5345 ( .A1(n7294), .A2(prog_data[5]), .B1(\mem[130][5] ), .B2(n7293), 
        .Z(n2578) );
  OA22D0 U5346 ( .A1(n7294), .A2(prog_data[4]), .B1(\mem[130][4] ), .B2(n7293), 
        .Z(n2577) );
  OA22D0 U5347 ( .A1(n7294), .A2(prog_data[3]), .B1(\mem[130][3] ), .B2(n7293), 
        .Z(n2576) );
  OA22D0 U5348 ( .A1(n7294), .A2(prog_data[2]), .B1(\mem[130][2] ), .B2(n7293), 
        .Z(n2575) );
  OA22D0 U5349 ( .A1(n7294), .A2(prog_data[1]), .B1(\mem[130][1] ), .B2(n7293), 
        .Z(n2574) );
  OA22D0 U5350 ( .A1(n7294), .A2(prog_data[0]), .B1(\mem[130][0] ), .B2(n7293), 
        .Z(n2573) );
  NR2D0 U5351 ( .A1(n7537), .A2(n7319), .ZN(n7295) );
  INVD0 U5352 ( .I(n7295), .ZN(n7296) );
  OA22D0 U5353 ( .A1(n7296), .A2(prog_data[15]), .B1(\mem[131][15] ), .B2(
        n7295), .Z(n2572) );
  OA22D0 U5354 ( .A1(n7296), .A2(prog_data[14]), .B1(\mem[131][14] ), .B2(
        n7295), .Z(n2571) );
  OA22D0 U5355 ( .A1(n7296), .A2(prog_data[13]), .B1(\mem[131][13] ), .B2(
        n7295), .Z(n2570) );
  OA22D0 U5356 ( .A1(n7296), .A2(prog_data[12]), .B1(\mem[131][12] ), .B2(
        n7295), .Z(n2569) );
  OA22D0 U5357 ( .A1(n7296), .A2(prog_data[11]), .B1(\mem[131][11] ), .B2(
        n7295), .Z(n2568) );
  OA22D0 U5358 ( .A1(n7296), .A2(prog_data[10]), .B1(\mem[131][10] ), .B2(
        n7295), .Z(n2567) );
  OA22D0 U5359 ( .A1(n7296), .A2(prog_data[9]), .B1(\mem[131][9] ), .B2(n7295), 
        .Z(n2566) );
  OA22D0 U5360 ( .A1(n7296), .A2(prog_data[8]), .B1(\mem[131][8] ), .B2(n7295), 
        .Z(n2565) );
  OA22D0 U5361 ( .A1(n7296), .A2(prog_data[7]), .B1(\mem[131][7] ), .B2(n7295), 
        .Z(n2564) );
  OA22D0 U5362 ( .A1(n7296), .A2(prog_data[6]), .B1(\mem[131][6] ), .B2(n7295), 
        .Z(n2563) );
  OA22D0 U5363 ( .A1(n7296), .A2(prog_data[5]), .B1(\mem[131][5] ), .B2(n7295), 
        .Z(n2562) );
  OA22D0 U5364 ( .A1(n7296), .A2(prog_data[4]), .B1(\mem[131][4] ), .B2(n7295), 
        .Z(n2561) );
  OA22D0 U5365 ( .A1(n7296), .A2(prog_data[3]), .B1(\mem[131][3] ), .B2(n7295), 
        .Z(n2560) );
  OA22D0 U5366 ( .A1(n7296), .A2(prog_data[2]), .B1(\mem[131][2] ), .B2(n7295), 
        .Z(n2559) );
  OA22D0 U5367 ( .A1(n7296), .A2(prog_data[1]), .B1(\mem[131][1] ), .B2(n7295), 
        .Z(n2558) );
  OA22D0 U5368 ( .A1(n7296), .A2(prog_data[0]), .B1(\mem[131][0] ), .B2(n7295), 
        .Z(n2557) );
  NR2D0 U5369 ( .A1(n7540), .A2(n7319), .ZN(n7297) );
  INVD0 U5370 ( .I(n7297), .ZN(n7298) );
  OA22D0 U5371 ( .A1(n7298), .A2(prog_data[15]), .B1(\mem[132][15] ), .B2(
        n7297), .Z(n2556) );
  OA22D0 U5372 ( .A1(n7298), .A2(prog_data[14]), .B1(\mem[132][14] ), .B2(
        n7297), .Z(n2555) );
  OA22D0 U5373 ( .A1(n7298), .A2(prog_data[13]), .B1(\mem[132][13] ), .B2(
        n7297), .Z(n2554) );
  OA22D0 U5374 ( .A1(n7298), .A2(prog_data[12]), .B1(\mem[132][12] ), .B2(
        n7297), .Z(n2553) );
  OA22D0 U5375 ( .A1(n7298), .A2(prog_data[11]), .B1(\mem[132][11] ), .B2(
        n7297), .Z(n2552) );
  OA22D0 U5376 ( .A1(n7298), .A2(prog_data[10]), .B1(\mem[132][10] ), .B2(
        n7297), .Z(n2551) );
  OA22D0 U5377 ( .A1(n7298), .A2(prog_data[9]), .B1(\mem[132][9] ), .B2(n7297), 
        .Z(n2550) );
  OA22D0 U5378 ( .A1(n7298), .A2(prog_data[8]), .B1(\mem[132][8] ), .B2(n7297), 
        .Z(n2549) );
  OA22D0 U5379 ( .A1(n7298), .A2(prog_data[7]), .B1(\mem[132][7] ), .B2(n7297), 
        .Z(n2548) );
  OA22D0 U5380 ( .A1(n7298), .A2(prog_data[6]), .B1(\mem[132][6] ), .B2(n7297), 
        .Z(n2547) );
  OA22D0 U5381 ( .A1(n7298), .A2(prog_data[5]), .B1(\mem[132][5] ), .B2(n7297), 
        .Z(n2546) );
  OA22D0 U5382 ( .A1(n7298), .A2(prog_data[4]), .B1(\mem[132][4] ), .B2(n7297), 
        .Z(n2545) );
  OA22D0 U5383 ( .A1(n7298), .A2(prog_data[3]), .B1(\mem[132][3] ), .B2(n7297), 
        .Z(n2544) );
  OA22D0 U5384 ( .A1(n7298), .A2(prog_data[2]), .B1(\mem[132][2] ), .B2(n7297), 
        .Z(n2543) );
  OA22D0 U5385 ( .A1(n7298), .A2(prog_data[1]), .B1(\mem[132][1] ), .B2(n7297), 
        .Z(n2542) );
  OA22D0 U5386 ( .A1(n7298), .A2(prog_data[0]), .B1(\mem[132][0] ), .B2(n7297), 
        .Z(n2541) );
  NR2D0 U5387 ( .A1(n7543), .A2(n7319), .ZN(n7299) );
  INVD0 U5388 ( .I(n7299), .ZN(n7300) );
  OA22D0 U5389 ( .A1(n7300), .A2(prog_data[15]), .B1(\mem[133][15] ), .B2(
        n7299), .Z(n2540) );
  OA22D0 U5390 ( .A1(n7300), .A2(prog_data[14]), .B1(\mem[133][14] ), .B2(
        n7299), .Z(n2539) );
  OA22D0 U5391 ( .A1(n7300), .A2(prog_data[13]), .B1(\mem[133][13] ), .B2(
        n7299), .Z(n2538) );
  OA22D0 U5392 ( .A1(n7300), .A2(prog_data[12]), .B1(\mem[133][12] ), .B2(
        n7299), .Z(n2537) );
  OA22D0 U5393 ( .A1(n7300), .A2(prog_data[11]), .B1(\mem[133][11] ), .B2(
        n7299), .Z(n2536) );
  OA22D0 U5394 ( .A1(n7300), .A2(prog_data[10]), .B1(\mem[133][10] ), .B2(
        n7299), .Z(n2535) );
  OA22D0 U5395 ( .A1(n7300), .A2(prog_data[9]), .B1(\mem[133][9] ), .B2(n7299), 
        .Z(n2534) );
  OA22D0 U5396 ( .A1(n7300), .A2(prog_data[8]), .B1(\mem[133][8] ), .B2(n7299), 
        .Z(n2533) );
  OA22D0 U5397 ( .A1(n7300), .A2(prog_data[7]), .B1(\mem[133][7] ), .B2(n7299), 
        .Z(n2532) );
  OA22D0 U5398 ( .A1(n7300), .A2(prog_data[6]), .B1(\mem[133][6] ), .B2(n7299), 
        .Z(n2531) );
  OA22D0 U5399 ( .A1(n7300), .A2(prog_data[5]), .B1(\mem[133][5] ), .B2(n7299), 
        .Z(n2530) );
  OA22D0 U5400 ( .A1(n7300), .A2(prog_data[4]), .B1(\mem[133][4] ), .B2(n7299), 
        .Z(n2529) );
  OA22D0 U5401 ( .A1(n7300), .A2(prog_data[3]), .B1(\mem[133][3] ), .B2(n7299), 
        .Z(n2528) );
  OA22D0 U5402 ( .A1(n7300), .A2(prog_data[2]), .B1(\mem[133][2] ), .B2(n7299), 
        .Z(n2527) );
  OA22D0 U5403 ( .A1(n7300), .A2(prog_data[1]), .B1(\mem[133][1] ), .B2(n7299), 
        .Z(n2526) );
  OA22D0 U5404 ( .A1(n7300), .A2(prog_data[0]), .B1(\mem[133][0] ), .B2(n7299), 
        .Z(n2525) );
  NR2D0 U5405 ( .A1(n7546), .A2(n7319), .ZN(n7301) );
  INVD0 U5406 ( .I(n7301), .ZN(n7302) );
  OA22D0 U5407 ( .A1(n7302), .A2(prog_data[15]), .B1(\mem[134][15] ), .B2(
        n7301), .Z(n2524) );
  OA22D0 U5408 ( .A1(n7302), .A2(prog_data[14]), .B1(\mem[134][14] ), .B2(
        n7301), .Z(n2523) );
  OA22D0 U5409 ( .A1(n7302), .A2(prog_data[13]), .B1(\mem[134][13] ), .B2(
        n7301), .Z(n2522) );
  OA22D0 U5410 ( .A1(n7302), .A2(prog_data[12]), .B1(\mem[134][12] ), .B2(
        n7301), .Z(n2521) );
  OA22D0 U5411 ( .A1(n7302), .A2(prog_data[11]), .B1(\mem[134][11] ), .B2(
        n7301), .Z(n2520) );
  OA22D0 U5412 ( .A1(n7302), .A2(prog_data[10]), .B1(\mem[134][10] ), .B2(
        n7301), .Z(n2519) );
  OA22D0 U5413 ( .A1(n7302), .A2(prog_data[9]), .B1(\mem[134][9] ), .B2(n7301), 
        .Z(n2518) );
  OA22D0 U5414 ( .A1(n7302), .A2(prog_data[8]), .B1(\mem[134][8] ), .B2(n7301), 
        .Z(n2517) );
  OA22D0 U5415 ( .A1(n7302), .A2(prog_data[7]), .B1(\mem[134][7] ), .B2(n7301), 
        .Z(n2516) );
  OA22D0 U5416 ( .A1(n7302), .A2(prog_data[6]), .B1(\mem[134][6] ), .B2(n7301), 
        .Z(n2515) );
  OA22D0 U5417 ( .A1(n7302), .A2(prog_data[5]), .B1(\mem[134][5] ), .B2(n7301), 
        .Z(n2514) );
  OA22D0 U5418 ( .A1(n7302), .A2(prog_data[4]), .B1(\mem[134][4] ), .B2(n7301), 
        .Z(n2513) );
  OA22D0 U5419 ( .A1(n7302), .A2(prog_data[3]), .B1(\mem[134][3] ), .B2(n7301), 
        .Z(n2512) );
  OA22D0 U5420 ( .A1(n7302), .A2(prog_data[2]), .B1(\mem[134][2] ), .B2(n7301), 
        .Z(n2511) );
  OA22D0 U5421 ( .A1(n7302), .A2(prog_data[1]), .B1(\mem[134][1] ), .B2(n7301), 
        .Z(n2510) );
  OA22D0 U5422 ( .A1(n7302), .A2(prog_data[0]), .B1(\mem[134][0] ), .B2(n7301), 
        .Z(n2509) );
  NR2D0 U5423 ( .A1(n7549), .A2(n7319), .ZN(n7303) );
  INVD0 U5424 ( .I(n7303), .ZN(n7304) );
  OA22D0 U5425 ( .A1(n7304), .A2(prog_data[15]), .B1(\mem[135][15] ), .B2(
        n7303), .Z(n2508) );
  OA22D0 U5426 ( .A1(n7304), .A2(prog_data[14]), .B1(\mem[135][14] ), .B2(
        n7303), .Z(n2507) );
  OA22D0 U5427 ( .A1(n7304), .A2(prog_data[13]), .B1(\mem[135][13] ), .B2(
        n7303), .Z(n2506) );
  OA22D0 U5428 ( .A1(n7304), .A2(prog_data[12]), .B1(\mem[135][12] ), .B2(
        n7303), .Z(n2505) );
  OA22D0 U5429 ( .A1(n7304), .A2(prog_data[11]), .B1(\mem[135][11] ), .B2(
        n7303), .Z(n2504) );
  OA22D0 U5430 ( .A1(n7304), .A2(prog_data[10]), .B1(\mem[135][10] ), .B2(
        n7303), .Z(n2503) );
  OA22D0 U5431 ( .A1(n7304), .A2(prog_data[9]), .B1(\mem[135][9] ), .B2(n7303), 
        .Z(n2502) );
  OA22D0 U5432 ( .A1(n7304), .A2(prog_data[8]), .B1(\mem[135][8] ), .B2(n7303), 
        .Z(n2501) );
  OA22D0 U5433 ( .A1(n7304), .A2(prog_data[7]), .B1(\mem[135][7] ), .B2(n7303), 
        .Z(n2500) );
  OA22D0 U5434 ( .A1(n7304), .A2(prog_data[6]), .B1(\mem[135][6] ), .B2(n7303), 
        .Z(n2499) );
  OA22D0 U5435 ( .A1(n7304), .A2(prog_data[5]), .B1(\mem[135][5] ), .B2(n7303), 
        .Z(n2498) );
  OA22D0 U5436 ( .A1(n7304), .A2(prog_data[4]), .B1(\mem[135][4] ), .B2(n7303), 
        .Z(n2497) );
  OA22D0 U5437 ( .A1(n7304), .A2(prog_data[3]), .B1(\mem[135][3] ), .B2(n7303), 
        .Z(n2496) );
  OA22D0 U5438 ( .A1(n7304), .A2(prog_data[2]), .B1(\mem[135][2] ), .B2(n7303), 
        .Z(n2495) );
  OA22D0 U5439 ( .A1(n7304), .A2(prog_data[1]), .B1(\mem[135][1] ), .B2(n7303), 
        .Z(n2494) );
  OA22D0 U5440 ( .A1(n7304), .A2(prog_data[0]), .B1(\mem[135][0] ), .B2(n7303), 
        .Z(n2493) );
  INVD0 U5441 ( .I(n7305), .ZN(n7306) );
  OA22D0 U5442 ( .A1(n7306), .A2(prog_data[15]), .B1(\mem[136][15] ), .B2(
        n7305), .Z(n2492) );
  OA22D0 U5443 ( .A1(n7306), .A2(prog_data[14]), .B1(\mem[136][14] ), .B2(
        n7305), .Z(n2491) );
  OA22D0 U5444 ( .A1(n7306), .A2(prog_data[13]), .B1(\mem[136][13] ), .B2(
        n7305), .Z(n2490) );
  OA22D0 U5445 ( .A1(n7306), .A2(prog_data[12]), .B1(\mem[136][12] ), .B2(
        n7305), .Z(n2489) );
  OA22D0 U5446 ( .A1(n7306), .A2(prog_data[11]), .B1(\mem[136][11] ), .B2(
        n7305), .Z(n2488) );
  OA22D0 U5447 ( .A1(n7306), .A2(prog_data[10]), .B1(\mem[136][10] ), .B2(
        n7305), .Z(n2487) );
  OA22D0 U5448 ( .A1(n7306), .A2(prog_data[9]), .B1(\mem[136][9] ), .B2(n7305), 
        .Z(n2486) );
  OA22D0 U5449 ( .A1(n7306), .A2(prog_data[8]), .B1(\mem[136][8] ), .B2(n7305), 
        .Z(n2485) );
  OA22D0 U5450 ( .A1(n7306), .A2(prog_data[7]), .B1(\mem[136][7] ), .B2(n7305), 
        .Z(n2484) );
  OA22D0 U5451 ( .A1(n7306), .A2(prog_data[6]), .B1(\mem[136][6] ), .B2(n7305), 
        .Z(n2483) );
  OA22D0 U5452 ( .A1(n7306), .A2(prog_data[5]), .B1(\mem[136][5] ), .B2(n7305), 
        .Z(n2482) );
  OA22D0 U5453 ( .A1(n7306), .A2(prog_data[4]), .B1(\mem[136][4] ), .B2(n7305), 
        .Z(n2481) );
  OA22D0 U5454 ( .A1(n7306), .A2(prog_data[3]), .B1(\mem[136][3] ), .B2(n7305), 
        .Z(n2480) );
  OA22D0 U5455 ( .A1(n7306), .A2(prog_data[2]), .B1(\mem[136][2] ), .B2(n7305), 
        .Z(n2479) );
  OA22D0 U5456 ( .A1(n7306), .A2(prog_data[1]), .B1(\mem[136][1] ), .B2(n7305), 
        .Z(n2478) );
  OA22D0 U5457 ( .A1(n7306), .A2(prog_data[0]), .B1(\mem[136][0] ), .B2(n7305), 
        .Z(n2477) );
  NR2D0 U5458 ( .A1(n7555), .A2(n7319), .ZN(n7307) );
  INVD0 U5459 ( .I(n7307), .ZN(n7308) );
  OA22D0 U5460 ( .A1(n7308), .A2(prog_data[15]), .B1(\mem[137][15] ), .B2(
        n7307), .Z(n2476) );
  OA22D0 U5461 ( .A1(n7308), .A2(prog_data[14]), .B1(\mem[137][14] ), .B2(
        n7307), .Z(n2475) );
  OA22D0 U5462 ( .A1(n7308), .A2(prog_data[13]), .B1(\mem[137][13] ), .B2(
        n7307), .Z(n2474) );
  OA22D0 U5463 ( .A1(n7308), .A2(prog_data[12]), .B1(\mem[137][12] ), .B2(
        n7307), .Z(n2473) );
  OA22D0 U5464 ( .A1(n7308), .A2(prog_data[11]), .B1(\mem[137][11] ), .B2(
        n7307), .Z(n2472) );
  OA22D0 U5465 ( .A1(n7308), .A2(prog_data[10]), .B1(\mem[137][10] ), .B2(
        n7307), .Z(n2471) );
  OA22D0 U5466 ( .A1(n7308), .A2(prog_data[9]), .B1(\mem[137][9] ), .B2(n7307), 
        .Z(n2470) );
  OA22D0 U5467 ( .A1(n7308), .A2(prog_data[8]), .B1(\mem[137][8] ), .B2(n7307), 
        .Z(n2469) );
  OA22D0 U5468 ( .A1(n7308), .A2(prog_data[7]), .B1(\mem[137][7] ), .B2(n7307), 
        .Z(n2468) );
  OA22D0 U5469 ( .A1(n7308), .A2(prog_data[6]), .B1(\mem[137][6] ), .B2(n7307), 
        .Z(n2467) );
  OA22D0 U5470 ( .A1(n7308), .A2(prog_data[5]), .B1(\mem[137][5] ), .B2(n7307), 
        .Z(n2466) );
  OA22D0 U5471 ( .A1(n7308), .A2(prog_data[4]), .B1(\mem[137][4] ), .B2(n7307), 
        .Z(n2465) );
  OA22D0 U5472 ( .A1(n7308), .A2(prog_data[3]), .B1(\mem[137][3] ), .B2(n7307), 
        .Z(n2464) );
  OA22D0 U5473 ( .A1(n7308), .A2(prog_data[2]), .B1(\mem[137][2] ), .B2(n7307), 
        .Z(n2463) );
  OA22D0 U5474 ( .A1(n7308), .A2(prog_data[1]), .B1(\mem[137][1] ), .B2(n7307), 
        .Z(n2462) );
  OA22D0 U5475 ( .A1(n7308), .A2(prog_data[0]), .B1(\mem[137][0] ), .B2(n7307), 
        .Z(n2461) );
  NR2D0 U5476 ( .A1(n7558), .A2(n7319), .ZN(n7309) );
  INVD0 U5477 ( .I(n7309), .ZN(n7310) );
  OA22D0 U5478 ( .A1(n7310), .A2(prog_data[15]), .B1(\mem[138][15] ), .B2(
        n7309), .Z(n2460) );
  OA22D0 U5479 ( .A1(n7310), .A2(prog_data[14]), .B1(\mem[138][14] ), .B2(
        n7309), .Z(n2459) );
  OA22D0 U5480 ( .A1(n7310), .A2(prog_data[13]), .B1(\mem[138][13] ), .B2(
        n7309), .Z(n2458) );
  OA22D0 U5481 ( .A1(n7310), .A2(prog_data[12]), .B1(\mem[138][12] ), .B2(
        n7309), .Z(n2457) );
  OA22D0 U5482 ( .A1(n7310), .A2(prog_data[11]), .B1(\mem[138][11] ), .B2(
        n7309), .Z(n2456) );
  OA22D0 U5483 ( .A1(n7310), .A2(prog_data[10]), .B1(\mem[138][10] ), .B2(
        n7309), .Z(n2455) );
  OA22D0 U5484 ( .A1(n7310), .A2(prog_data[9]), .B1(\mem[138][9] ), .B2(n7309), 
        .Z(n2454) );
  OA22D0 U5485 ( .A1(n7310), .A2(prog_data[8]), .B1(\mem[138][8] ), .B2(n7309), 
        .Z(n2453) );
  OA22D0 U5486 ( .A1(n7310), .A2(prog_data[7]), .B1(\mem[138][7] ), .B2(n7309), 
        .Z(n2452) );
  OA22D0 U5487 ( .A1(n7310), .A2(prog_data[6]), .B1(\mem[138][6] ), .B2(n7309), 
        .Z(n2451) );
  OA22D0 U5488 ( .A1(n7310), .A2(prog_data[5]), .B1(\mem[138][5] ), .B2(n7309), 
        .Z(n2450) );
  OA22D0 U5489 ( .A1(n7310), .A2(prog_data[4]), .B1(\mem[138][4] ), .B2(n7309), 
        .Z(n2449) );
  OA22D0 U5490 ( .A1(n7310), .A2(prog_data[3]), .B1(\mem[138][3] ), .B2(n7309), 
        .Z(n2448) );
  OA22D0 U5491 ( .A1(n7310), .A2(prog_data[2]), .B1(\mem[138][2] ), .B2(n7309), 
        .Z(n2447) );
  OA22D0 U5492 ( .A1(n7310), .A2(prog_data[1]), .B1(\mem[138][1] ), .B2(n7309), 
        .Z(n2446) );
  OA22D0 U5493 ( .A1(n7310), .A2(prog_data[0]), .B1(\mem[138][0] ), .B2(n7309), 
        .Z(n2445) );
  NR2D0 U5494 ( .A1(n7561), .A2(n7319), .ZN(n7311) );
  INVD0 U5495 ( .I(n7311), .ZN(n7312) );
  OA22D0 U5496 ( .A1(n7312), .A2(prog_data[15]), .B1(\mem[139][15] ), .B2(
        n7311), .Z(n2444) );
  OA22D0 U5497 ( .A1(n7312), .A2(prog_data[14]), .B1(\mem[139][14] ), .B2(
        n7311), .Z(n2443) );
  OA22D0 U5498 ( .A1(n7312), .A2(prog_data[13]), .B1(\mem[139][13] ), .B2(
        n7311), .Z(n2442) );
  OA22D0 U5499 ( .A1(n7312), .A2(prog_data[12]), .B1(\mem[139][12] ), .B2(
        n7311), .Z(n2441) );
  OA22D0 U5500 ( .A1(n7312), .A2(prog_data[11]), .B1(\mem[139][11] ), .B2(
        n7311), .Z(n2440) );
  OA22D0 U5501 ( .A1(n7312), .A2(prog_data[10]), .B1(\mem[139][10] ), .B2(
        n7311), .Z(n2439) );
  OA22D0 U5502 ( .A1(n7312), .A2(prog_data[9]), .B1(\mem[139][9] ), .B2(n7311), 
        .Z(n2438) );
  OA22D0 U5503 ( .A1(n7312), .A2(prog_data[8]), .B1(\mem[139][8] ), .B2(n7311), 
        .Z(n2437) );
  OA22D0 U5504 ( .A1(n7312), .A2(prog_data[7]), .B1(\mem[139][7] ), .B2(n7311), 
        .Z(n2436) );
  OA22D0 U5505 ( .A1(n7312), .A2(prog_data[6]), .B1(\mem[139][6] ), .B2(n7311), 
        .Z(n2435) );
  OA22D0 U5506 ( .A1(n7312), .A2(prog_data[5]), .B1(\mem[139][5] ), .B2(n7311), 
        .Z(n2434) );
  OA22D0 U5507 ( .A1(n7312), .A2(prog_data[4]), .B1(\mem[139][4] ), .B2(n7311), 
        .Z(n2433) );
  OA22D0 U5508 ( .A1(n7312), .A2(prog_data[3]), .B1(\mem[139][3] ), .B2(n7311), 
        .Z(n2432) );
  OA22D0 U5509 ( .A1(n7312), .A2(prog_data[2]), .B1(\mem[139][2] ), .B2(n7311), 
        .Z(n2431) );
  OA22D0 U5510 ( .A1(n7312), .A2(prog_data[1]), .B1(\mem[139][1] ), .B2(n7311), 
        .Z(n2430) );
  OA22D0 U5511 ( .A1(n7312), .A2(prog_data[0]), .B1(\mem[139][0] ), .B2(n7311), 
        .Z(n2429) );
  NR2D0 U5512 ( .A1(n7564), .A2(n7319), .ZN(n7313) );
  INVD0 U5513 ( .I(n7313), .ZN(n7314) );
  OA22D0 U5514 ( .A1(n7314), .A2(prog_data[15]), .B1(\mem[140][15] ), .B2(
        n7313), .Z(n2428) );
  OA22D0 U5515 ( .A1(n7314), .A2(prog_data[14]), .B1(\mem[140][14] ), .B2(
        n7313), .Z(n2427) );
  OA22D0 U5516 ( .A1(n7314), .A2(prog_data[13]), .B1(\mem[140][13] ), .B2(
        n7313), .Z(n2426) );
  OA22D0 U5517 ( .A1(n7314), .A2(prog_data[12]), .B1(\mem[140][12] ), .B2(
        n7313), .Z(n2425) );
  OA22D0 U5518 ( .A1(n7314), .A2(prog_data[11]), .B1(\mem[140][11] ), .B2(
        n7313), .Z(n2424) );
  OA22D0 U5519 ( .A1(n7314), .A2(prog_data[10]), .B1(\mem[140][10] ), .B2(
        n7313), .Z(n2423) );
  OA22D0 U5520 ( .A1(n7314), .A2(prog_data[9]), .B1(\mem[140][9] ), .B2(n7313), 
        .Z(n2422) );
  OA22D0 U5521 ( .A1(n7314), .A2(prog_data[8]), .B1(\mem[140][8] ), .B2(n7313), 
        .Z(n2421) );
  OA22D0 U5522 ( .A1(n7314), .A2(prog_data[7]), .B1(\mem[140][7] ), .B2(n7313), 
        .Z(n2420) );
  OA22D0 U5523 ( .A1(n7314), .A2(prog_data[6]), .B1(\mem[140][6] ), .B2(n7313), 
        .Z(n2419) );
  OA22D0 U5524 ( .A1(n7314), .A2(prog_data[5]), .B1(\mem[140][5] ), .B2(n7313), 
        .Z(n2418) );
  OA22D0 U5525 ( .A1(n7314), .A2(prog_data[4]), .B1(\mem[140][4] ), .B2(n7313), 
        .Z(n2417) );
  OA22D0 U5526 ( .A1(n7314), .A2(prog_data[3]), .B1(\mem[140][3] ), .B2(n7313), 
        .Z(n2416) );
  OA22D0 U5527 ( .A1(n7314), .A2(prog_data[2]), .B1(\mem[140][2] ), .B2(n7313), 
        .Z(n2415) );
  OA22D0 U5528 ( .A1(n7314), .A2(prog_data[1]), .B1(\mem[140][1] ), .B2(n7313), 
        .Z(n2414) );
  OA22D0 U5529 ( .A1(n7314), .A2(prog_data[0]), .B1(\mem[140][0] ), .B2(n7313), 
        .Z(n2413) );
  NR2D0 U5530 ( .A1(n7567), .A2(n7319), .ZN(n7315) );
  INVD0 U5531 ( .I(n7315), .ZN(n7316) );
  OA22D0 U5532 ( .A1(n7316), .A2(prog_data[15]), .B1(\mem[141][15] ), .B2(
        n7315), .Z(n2412) );
  OA22D0 U5533 ( .A1(n7316), .A2(prog_data[14]), .B1(\mem[141][14] ), .B2(
        n7315), .Z(n2411) );
  OA22D0 U5534 ( .A1(n7316), .A2(prog_data[13]), .B1(\mem[141][13] ), .B2(
        n7315), .Z(n2410) );
  OA22D0 U5535 ( .A1(n7316), .A2(prog_data[12]), .B1(\mem[141][12] ), .B2(
        n7315), .Z(n2409) );
  OA22D0 U5536 ( .A1(n7316), .A2(prog_data[11]), .B1(\mem[141][11] ), .B2(
        n7315), .Z(n2408) );
  OA22D0 U5537 ( .A1(n7316), .A2(prog_data[10]), .B1(\mem[141][10] ), .B2(
        n7315), .Z(n2407) );
  OA22D0 U5538 ( .A1(n7316), .A2(prog_data[9]), .B1(\mem[141][9] ), .B2(n7315), 
        .Z(n2406) );
  OA22D0 U5539 ( .A1(n7316), .A2(prog_data[8]), .B1(\mem[141][8] ), .B2(n7315), 
        .Z(n2405) );
  OA22D0 U5540 ( .A1(n7316), .A2(prog_data[7]), .B1(\mem[141][7] ), .B2(n7315), 
        .Z(n2404) );
  OA22D0 U5541 ( .A1(n7316), .A2(prog_data[6]), .B1(\mem[141][6] ), .B2(n7315), 
        .Z(n2403) );
  OA22D0 U5542 ( .A1(n7316), .A2(prog_data[5]), .B1(\mem[141][5] ), .B2(n7315), 
        .Z(n2402) );
  OA22D0 U5543 ( .A1(n7316), .A2(prog_data[4]), .B1(\mem[141][4] ), .B2(n7315), 
        .Z(n2401) );
  OA22D0 U5544 ( .A1(n7316), .A2(prog_data[3]), .B1(\mem[141][3] ), .B2(n7315), 
        .Z(n2400) );
  OA22D0 U5545 ( .A1(n7316), .A2(prog_data[2]), .B1(\mem[141][2] ), .B2(n7315), 
        .Z(n2399) );
  OA22D0 U5546 ( .A1(n7316), .A2(prog_data[1]), .B1(\mem[141][1] ), .B2(n7315), 
        .Z(n2398) );
  OA22D0 U5547 ( .A1(n7316), .A2(prog_data[0]), .B1(\mem[141][0] ), .B2(n7315), 
        .Z(n2397) );
  NR2D0 U5548 ( .A1(n7570), .A2(n7319), .ZN(n7317) );
  INVD0 U5549 ( .I(n7317), .ZN(n7318) );
  OA22D0 U5550 ( .A1(n7318), .A2(prog_data[15]), .B1(\mem[142][15] ), .B2(
        n7317), .Z(n2396) );
  OA22D0 U5551 ( .A1(n7318), .A2(prog_data[14]), .B1(\mem[142][14] ), .B2(
        n7317), .Z(n2395) );
  OA22D0 U5552 ( .A1(n7318), .A2(prog_data[13]), .B1(\mem[142][13] ), .B2(
        n7317), .Z(n2394) );
  OA22D0 U5553 ( .A1(n7318), .A2(prog_data[12]), .B1(\mem[142][12] ), .B2(
        n7317), .Z(n2393) );
  OA22D0 U5554 ( .A1(n7318), .A2(prog_data[11]), .B1(\mem[142][11] ), .B2(
        n7317), .Z(n2392) );
  OA22D0 U5555 ( .A1(n7318), .A2(prog_data[10]), .B1(\mem[142][10] ), .B2(
        n7317), .Z(n2391) );
  OA22D0 U5556 ( .A1(n7318), .A2(prog_data[9]), .B1(\mem[142][9] ), .B2(n7317), 
        .Z(n2390) );
  OA22D0 U5557 ( .A1(n7318), .A2(prog_data[8]), .B1(\mem[142][8] ), .B2(n7317), 
        .Z(n2389) );
  OA22D0 U5558 ( .A1(n7318), .A2(prog_data[7]), .B1(\mem[142][7] ), .B2(n7317), 
        .Z(n2388) );
  OA22D0 U5559 ( .A1(n7318), .A2(prog_data[6]), .B1(\mem[142][6] ), .B2(n7317), 
        .Z(n2387) );
  OA22D0 U5560 ( .A1(n7318), .A2(prog_data[5]), .B1(\mem[142][5] ), .B2(n7317), 
        .Z(n2386) );
  OA22D0 U5561 ( .A1(n7318), .A2(prog_data[4]), .B1(\mem[142][4] ), .B2(n7317), 
        .Z(n2385) );
  OA22D0 U5562 ( .A1(n7318), .A2(prog_data[3]), .B1(\mem[142][3] ), .B2(n7317), 
        .Z(n2384) );
  OA22D0 U5563 ( .A1(n7318), .A2(prog_data[2]), .B1(\mem[142][2] ), .B2(n7317), 
        .Z(n2383) );
  OA22D0 U5564 ( .A1(n7318), .A2(prog_data[1]), .B1(\mem[142][1] ), .B2(n7317), 
        .Z(n2382) );
  OA22D0 U5565 ( .A1(n7318), .A2(prog_data[0]), .B1(\mem[142][0] ), .B2(n7317), 
        .Z(n2381) );
  NR2D0 U5566 ( .A1(n7574), .A2(n7319), .ZN(n7320) );
  INVD0 U5567 ( .I(n7320), .ZN(n7321) );
  OA22D0 U5568 ( .A1(n7321), .A2(prog_data[15]), .B1(\mem[143][15] ), .B2(
        n7320), .Z(n2380) );
  OA22D0 U5569 ( .A1(n7321), .A2(prog_data[14]), .B1(\mem[143][14] ), .B2(
        n7320), .Z(n2379) );
  OA22D0 U5570 ( .A1(n7321), .A2(prog_data[13]), .B1(\mem[143][13] ), .B2(
        n7320), .Z(n2378) );
  OA22D0 U5571 ( .A1(n7321), .A2(prog_data[12]), .B1(\mem[143][12] ), .B2(
        n7320), .Z(n2377) );
  OA22D0 U5572 ( .A1(n7321), .A2(prog_data[11]), .B1(\mem[143][11] ), .B2(
        n7320), .Z(n2376) );
  OA22D0 U5573 ( .A1(n7321), .A2(prog_data[10]), .B1(\mem[143][10] ), .B2(
        n7320), .Z(n2375) );
  OA22D0 U5574 ( .A1(n7321), .A2(prog_data[9]), .B1(\mem[143][9] ), .B2(n7320), 
        .Z(n2374) );
  OA22D0 U5575 ( .A1(n7321), .A2(prog_data[8]), .B1(\mem[143][8] ), .B2(n7320), 
        .Z(n2373) );
  OA22D0 U5576 ( .A1(n7321), .A2(prog_data[7]), .B1(\mem[143][7] ), .B2(n7320), 
        .Z(n2372) );
  OA22D0 U5577 ( .A1(n7321), .A2(prog_data[6]), .B1(\mem[143][6] ), .B2(n7320), 
        .Z(n2371) );
  OA22D0 U5578 ( .A1(n7321), .A2(prog_data[5]), .B1(\mem[143][5] ), .B2(n7320), 
        .Z(n2370) );
  OA22D0 U5579 ( .A1(n7321), .A2(prog_data[4]), .B1(\mem[143][4] ), .B2(n7320), 
        .Z(n2369) );
  OA22D0 U5580 ( .A1(n7321), .A2(prog_data[3]), .B1(\mem[143][3] ), .B2(n7320), 
        .Z(n2368) );
  OA22D0 U5581 ( .A1(n7321), .A2(prog_data[2]), .B1(\mem[143][2] ), .B2(n7320), 
        .Z(n2367) );
  OA22D0 U5582 ( .A1(n7321), .A2(prog_data[1]), .B1(\mem[143][1] ), .B2(n7320), 
        .Z(n2366) );
  OA22D0 U5583 ( .A1(n7321), .A2(prog_data[0]), .B1(\mem[143][0] ), .B2(n7320), 
        .Z(n2365) );
  NR2D0 U5584 ( .A1(n7323), .A2(n7322), .ZN(n7526) );
  CKND2D0 U5585 ( .A1(n7324), .A2(n7526), .ZN(n7355) );
  NR2D0 U5586 ( .A1(n7528), .A2(n7355), .ZN(n7325) );
  OA22D0 U5587 ( .A1(n7326), .A2(prog_data[15]), .B1(\mem[144][15] ), .B2(
        n7325), .Z(n2364) );
  OA22D0 U5588 ( .A1(n7326), .A2(prog_data[14]), .B1(\mem[144][14] ), .B2(
        n7325), .Z(n2363) );
  OA22D0 U5589 ( .A1(n7326), .A2(prog_data[13]), .B1(\mem[144][13] ), .B2(
        n7325), .Z(n2362) );
  OA22D0 U5590 ( .A1(n7326), .A2(prog_data[12]), .B1(\mem[144][12] ), .B2(
        n7325), .Z(n2361) );
  OA22D0 U5591 ( .A1(n7326), .A2(prog_data[11]), .B1(\mem[144][11] ), .B2(
        n7325), .Z(n2360) );
  OA22D0 U5592 ( .A1(n7326), .A2(prog_data[10]), .B1(\mem[144][10] ), .B2(
        n7325), .Z(n2359) );
  OA22D0 U5593 ( .A1(n7326), .A2(prog_data[9]), .B1(\mem[144][9] ), .B2(n7325), 
        .Z(n2358) );
  OA22D0 U5594 ( .A1(n7326), .A2(prog_data[8]), .B1(\mem[144][8] ), .B2(n7325), 
        .Z(n2357) );
  OA22D0 U5595 ( .A1(n7326), .A2(prog_data[7]), .B1(\mem[144][7] ), .B2(n7325), 
        .Z(n2356) );
  OA22D0 U5596 ( .A1(n7326), .A2(prog_data[6]), .B1(\mem[144][6] ), .B2(n7325), 
        .Z(n2355) );
  OA22D0 U5597 ( .A1(n7326), .A2(prog_data[5]), .B1(\mem[144][5] ), .B2(n7325), 
        .Z(n2354) );
  OA22D0 U5598 ( .A1(n7326), .A2(prog_data[4]), .B1(\mem[144][4] ), .B2(n7325), 
        .Z(n2353) );
  OA22D0 U5599 ( .A1(n7326), .A2(prog_data[3]), .B1(\mem[144][3] ), .B2(n7325), 
        .Z(n2352) );
  OA22D0 U5600 ( .A1(n7326), .A2(prog_data[2]), .B1(\mem[144][2] ), .B2(n7325), 
        .Z(n2351) );
  OA22D0 U5601 ( .A1(n7326), .A2(prog_data[1]), .B1(\mem[144][1] ), .B2(n7325), 
        .Z(n2350) );
  OA22D0 U5602 ( .A1(n7326), .A2(prog_data[0]), .B1(\mem[144][0] ), .B2(n7325), 
        .Z(n2349) );
  NR2D0 U5603 ( .A1(n7531), .A2(n7355), .ZN(n7327) );
  INVD0 U5604 ( .I(n7327), .ZN(n7328) );
  OA22D0 U5605 ( .A1(n7328), .A2(prog_data[15]), .B1(\mem[145][15] ), .B2(
        n7327), .Z(n2348) );
  OA22D0 U5606 ( .A1(n7328), .A2(prog_data[14]), .B1(\mem[145][14] ), .B2(
        n7327), .Z(n2347) );
  OA22D0 U5607 ( .A1(n7328), .A2(prog_data[13]), .B1(\mem[145][13] ), .B2(
        n7327), .Z(n2346) );
  OA22D0 U5608 ( .A1(n7328), .A2(prog_data[12]), .B1(\mem[145][12] ), .B2(
        n7327), .Z(n2345) );
  OA22D0 U5609 ( .A1(n7328), .A2(prog_data[11]), .B1(\mem[145][11] ), .B2(
        n7327), .Z(n2344) );
  OA22D0 U5610 ( .A1(n7328), .A2(prog_data[10]), .B1(\mem[145][10] ), .B2(
        n7327), .Z(n2343) );
  OA22D0 U5611 ( .A1(n7328), .A2(prog_data[9]), .B1(\mem[145][9] ), .B2(n7327), 
        .Z(n2342) );
  OA22D0 U5612 ( .A1(n7328), .A2(prog_data[8]), .B1(\mem[145][8] ), .B2(n7327), 
        .Z(n2341) );
  OA22D0 U5613 ( .A1(n7328), .A2(prog_data[7]), .B1(\mem[145][7] ), .B2(n7327), 
        .Z(n2340) );
  OA22D0 U5614 ( .A1(n7328), .A2(prog_data[6]), .B1(\mem[145][6] ), .B2(n7327), 
        .Z(n2339) );
  OA22D0 U5615 ( .A1(n7328), .A2(prog_data[5]), .B1(\mem[145][5] ), .B2(n7327), 
        .Z(n2338) );
  OA22D0 U5616 ( .A1(n7328), .A2(prog_data[4]), .B1(\mem[145][4] ), .B2(n7327), 
        .Z(n2337) );
  OA22D0 U5617 ( .A1(n7328), .A2(prog_data[3]), .B1(\mem[145][3] ), .B2(n7327), 
        .Z(n2336) );
  OA22D0 U5618 ( .A1(n7328), .A2(prog_data[2]), .B1(\mem[145][2] ), .B2(n7327), 
        .Z(n2335) );
  OA22D0 U5619 ( .A1(n7328), .A2(prog_data[1]), .B1(\mem[145][1] ), .B2(n7327), 
        .Z(n2334) );
  OA22D0 U5620 ( .A1(n7328), .A2(prog_data[0]), .B1(\mem[145][0] ), .B2(n7327), 
        .Z(n2333) );
  NR2D0 U5621 ( .A1(n7534), .A2(n7355), .ZN(n7329) );
  INVD0 U5622 ( .I(n7329), .ZN(n7330) );
  OA22D0 U5623 ( .A1(n7330), .A2(prog_data[15]), .B1(\mem[146][15] ), .B2(
        n7329), .Z(n2332) );
  OA22D0 U5624 ( .A1(n7330), .A2(prog_data[14]), .B1(\mem[146][14] ), .B2(
        n7329), .Z(n2331) );
  OA22D0 U5625 ( .A1(n7330), .A2(prog_data[13]), .B1(\mem[146][13] ), .B2(
        n7329), .Z(n2330) );
  OA22D0 U5626 ( .A1(n7330), .A2(prog_data[12]), .B1(\mem[146][12] ), .B2(
        n7329), .Z(n2329) );
  OA22D0 U5627 ( .A1(n7330), .A2(prog_data[11]), .B1(\mem[146][11] ), .B2(
        n7329), .Z(n2328) );
  OA22D0 U5628 ( .A1(n7330), .A2(prog_data[10]), .B1(\mem[146][10] ), .B2(
        n7329), .Z(n2327) );
  OA22D0 U5629 ( .A1(n7330), .A2(prog_data[9]), .B1(\mem[146][9] ), .B2(n7329), 
        .Z(n2326) );
  OA22D0 U5630 ( .A1(n7330), .A2(prog_data[8]), .B1(\mem[146][8] ), .B2(n7329), 
        .Z(n2325) );
  OA22D0 U5631 ( .A1(n7330), .A2(prog_data[7]), .B1(\mem[146][7] ), .B2(n7329), 
        .Z(n2324) );
  OA22D0 U5632 ( .A1(n7330), .A2(prog_data[6]), .B1(\mem[146][6] ), .B2(n7329), 
        .Z(n2323) );
  OA22D0 U5633 ( .A1(n7330), .A2(prog_data[5]), .B1(\mem[146][5] ), .B2(n7329), 
        .Z(n2322) );
  OA22D0 U5634 ( .A1(n7330), .A2(prog_data[4]), .B1(\mem[146][4] ), .B2(n7329), 
        .Z(n2321) );
  OA22D0 U5635 ( .A1(n7330), .A2(prog_data[3]), .B1(\mem[146][3] ), .B2(n7329), 
        .Z(n2320) );
  OA22D0 U5636 ( .A1(n7330), .A2(prog_data[2]), .B1(\mem[146][2] ), .B2(n7329), 
        .Z(n2319) );
  OA22D0 U5637 ( .A1(n7330), .A2(prog_data[1]), .B1(\mem[146][1] ), .B2(n7329), 
        .Z(n2318) );
  OA22D0 U5638 ( .A1(n7330), .A2(prog_data[0]), .B1(\mem[146][0] ), .B2(n7329), 
        .Z(n2317) );
  NR2D0 U5639 ( .A1(n7537), .A2(n7355), .ZN(n7331) );
  INVD0 U5640 ( .I(n7331), .ZN(n7332) );
  OA22D0 U5641 ( .A1(n7332), .A2(prog_data[15]), .B1(\mem[147][15] ), .B2(
        n7331), .Z(n2316) );
  OA22D0 U5642 ( .A1(n7332), .A2(prog_data[14]), .B1(\mem[147][14] ), .B2(
        n7331), .Z(n2315) );
  OA22D0 U5643 ( .A1(n7332), .A2(prog_data[13]), .B1(\mem[147][13] ), .B2(
        n7331), .Z(n2314) );
  OA22D0 U5644 ( .A1(n7332), .A2(prog_data[12]), .B1(\mem[147][12] ), .B2(
        n7331), .Z(n2313) );
  OA22D0 U5645 ( .A1(n7332), .A2(prog_data[11]), .B1(\mem[147][11] ), .B2(
        n7331), .Z(n2312) );
  OA22D0 U5646 ( .A1(n7332), .A2(prog_data[10]), .B1(\mem[147][10] ), .B2(
        n7331), .Z(n2311) );
  OA22D0 U5647 ( .A1(n7332), .A2(prog_data[9]), .B1(\mem[147][9] ), .B2(n7331), 
        .Z(n2310) );
  OA22D0 U5648 ( .A1(n7332), .A2(prog_data[8]), .B1(\mem[147][8] ), .B2(n7331), 
        .Z(n2309) );
  OA22D0 U5649 ( .A1(n7332), .A2(prog_data[7]), .B1(\mem[147][7] ), .B2(n7331), 
        .Z(n2308) );
  OA22D0 U5650 ( .A1(n7332), .A2(prog_data[6]), .B1(\mem[147][6] ), .B2(n7331), 
        .Z(n2307) );
  OA22D0 U5651 ( .A1(n7332), .A2(prog_data[5]), .B1(\mem[147][5] ), .B2(n7331), 
        .Z(n2306) );
  OA22D0 U5652 ( .A1(n7332), .A2(prog_data[4]), .B1(\mem[147][4] ), .B2(n7331), 
        .Z(n2305) );
  OA22D0 U5653 ( .A1(n7332), .A2(prog_data[3]), .B1(\mem[147][3] ), .B2(n7331), 
        .Z(n2304) );
  OA22D0 U5654 ( .A1(n7332), .A2(prog_data[2]), .B1(\mem[147][2] ), .B2(n7331), 
        .Z(n2303) );
  OA22D0 U5655 ( .A1(n7332), .A2(prog_data[1]), .B1(\mem[147][1] ), .B2(n7331), 
        .Z(n2302) );
  OA22D0 U5656 ( .A1(n7332), .A2(prog_data[0]), .B1(\mem[147][0] ), .B2(n7331), 
        .Z(n2301) );
  NR2D0 U5657 ( .A1(n7540), .A2(n7355), .ZN(n7333) );
  INVD0 U5658 ( .I(n7333), .ZN(n7334) );
  OA22D0 U5659 ( .A1(n7334), .A2(prog_data[15]), .B1(\mem[148][15] ), .B2(
        n7333), .Z(n2300) );
  OA22D0 U5660 ( .A1(n7334), .A2(prog_data[14]), .B1(\mem[148][14] ), .B2(
        n7333), .Z(n2299) );
  OA22D0 U5661 ( .A1(n7334), .A2(prog_data[13]), .B1(\mem[148][13] ), .B2(
        n7333), .Z(n2298) );
  OA22D0 U5662 ( .A1(n7334), .A2(prog_data[12]), .B1(\mem[148][12] ), .B2(
        n7333), .Z(n2297) );
  OA22D0 U5663 ( .A1(n7334), .A2(prog_data[11]), .B1(\mem[148][11] ), .B2(
        n7333), .Z(n2296) );
  OA22D0 U5664 ( .A1(n7334), .A2(prog_data[10]), .B1(\mem[148][10] ), .B2(
        n7333), .Z(n2295) );
  OA22D0 U5665 ( .A1(n7334), .A2(prog_data[9]), .B1(\mem[148][9] ), .B2(n7333), 
        .Z(n2294) );
  OA22D0 U5666 ( .A1(n7334), .A2(prog_data[8]), .B1(\mem[148][8] ), .B2(n7333), 
        .Z(n2293) );
  OA22D0 U5667 ( .A1(n7334), .A2(prog_data[7]), .B1(\mem[148][7] ), .B2(n7333), 
        .Z(n2292) );
  OA22D0 U5668 ( .A1(n7334), .A2(prog_data[6]), .B1(\mem[148][6] ), .B2(n7333), 
        .Z(n2291) );
  OA22D0 U5669 ( .A1(n7334), .A2(prog_data[5]), .B1(\mem[148][5] ), .B2(n7333), 
        .Z(n2290) );
  OA22D0 U5670 ( .A1(n7334), .A2(prog_data[4]), .B1(\mem[148][4] ), .B2(n7333), 
        .Z(n2289) );
  OA22D0 U5671 ( .A1(n7334), .A2(prog_data[3]), .B1(\mem[148][3] ), .B2(n7333), 
        .Z(n2288) );
  OA22D0 U5672 ( .A1(n7334), .A2(prog_data[2]), .B1(\mem[148][2] ), .B2(n7333), 
        .Z(n2287) );
  OA22D0 U5673 ( .A1(n7334), .A2(prog_data[1]), .B1(\mem[148][1] ), .B2(n7333), 
        .Z(n2286) );
  OA22D0 U5674 ( .A1(n7334), .A2(prog_data[0]), .B1(\mem[148][0] ), .B2(n7333), 
        .Z(n2285) );
  NR2D0 U5675 ( .A1(n7543), .A2(n7355), .ZN(n7335) );
  INVD0 U5676 ( .I(n7335), .ZN(n7336) );
  OA22D0 U5677 ( .A1(n7336), .A2(prog_data[15]), .B1(\mem[149][15] ), .B2(
        n7335), .Z(n2284) );
  OA22D0 U5678 ( .A1(n7336), .A2(prog_data[14]), .B1(\mem[149][14] ), .B2(
        n7335), .Z(n2283) );
  OA22D0 U5679 ( .A1(n7336), .A2(prog_data[13]), .B1(\mem[149][13] ), .B2(
        n7335), .Z(n2282) );
  OA22D0 U5680 ( .A1(n7336), .A2(prog_data[12]), .B1(\mem[149][12] ), .B2(
        n7335), .Z(n2281) );
  OA22D0 U5681 ( .A1(n7336), .A2(prog_data[11]), .B1(\mem[149][11] ), .B2(
        n7335), .Z(n2280) );
  OA22D0 U5682 ( .A1(n7336), .A2(prog_data[10]), .B1(\mem[149][10] ), .B2(
        n7335), .Z(n2279) );
  OA22D0 U5683 ( .A1(n7336), .A2(prog_data[9]), .B1(\mem[149][9] ), .B2(n7335), 
        .Z(n2278) );
  OA22D0 U5684 ( .A1(n7336), .A2(prog_data[8]), .B1(\mem[149][8] ), .B2(n7335), 
        .Z(n2277) );
  OA22D0 U5685 ( .A1(n7336), .A2(prog_data[7]), .B1(\mem[149][7] ), .B2(n7335), 
        .Z(n2276) );
  OA22D0 U5686 ( .A1(n7336), .A2(prog_data[6]), .B1(\mem[149][6] ), .B2(n7335), 
        .Z(n2275) );
  OA22D0 U5687 ( .A1(n7336), .A2(prog_data[5]), .B1(\mem[149][5] ), .B2(n7335), 
        .Z(n2274) );
  OA22D0 U5688 ( .A1(n7336), .A2(prog_data[4]), .B1(\mem[149][4] ), .B2(n7335), 
        .Z(n2273) );
  OA22D0 U5689 ( .A1(n7336), .A2(prog_data[3]), .B1(\mem[149][3] ), .B2(n7335), 
        .Z(n2272) );
  OA22D0 U5690 ( .A1(n7336), .A2(prog_data[2]), .B1(\mem[149][2] ), .B2(n7335), 
        .Z(n2271) );
  OA22D0 U5691 ( .A1(n7336), .A2(prog_data[1]), .B1(\mem[149][1] ), .B2(n7335), 
        .Z(n2270) );
  OA22D0 U5692 ( .A1(n7336), .A2(prog_data[0]), .B1(\mem[149][0] ), .B2(n7335), 
        .Z(n2269) );
  NR2D0 U5693 ( .A1(n7546), .A2(n7355), .ZN(n7337) );
  INVD0 U5694 ( .I(n7337), .ZN(n7338) );
  OA22D0 U5695 ( .A1(n7338), .A2(prog_data[15]), .B1(\mem[150][15] ), .B2(
        n7337), .Z(n2268) );
  OA22D0 U5696 ( .A1(n7338), .A2(prog_data[14]), .B1(\mem[150][14] ), .B2(
        n7337), .Z(n2267) );
  OA22D0 U5697 ( .A1(n7338), .A2(prog_data[13]), .B1(\mem[150][13] ), .B2(
        n7337), .Z(n2266) );
  OA22D0 U5698 ( .A1(n7338), .A2(prog_data[12]), .B1(\mem[150][12] ), .B2(
        n7337), .Z(n2265) );
  OA22D0 U5699 ( .A1(n7338), .A2(prog_data[11]), .B1(\mem[150][11] ), .B2(
        n7337), .Z(n2264) );
  OA22D0 U5700 ( .A1(n7338), .A2(prog_data[10]), .B1(\mem[150][10] ), .B2(
        n7337), .Z(n2263) );
  OA22D0 U5701 ( .A1(n7338), .A2(prog_data[9]), .B1(\mem[150][9] ), .B2(n7337), 
        .Z(n2262) );
  OA22D0 U5702 ( .A1(n7338), .A2(prog_data[8]), .B1(\mem[150][8] ), .B2(n7337), 
        .Z(n2261) );
  OA22D0 U5703 ( .A1(n7338), .A2(prog_data[7]), .B1(\mem[150][7] ), .B2(n7337), 
        .Z(n2260) );
  OA22D0 U5704 ( .A1(n7338), .A2(prog_data[6]), .B1(\mem[150][6] ), .B2(n7337), 
        .Z(n2259) );
  OA22D0 U5705 ( .A1(n7338), .A2(prog_data[5]), .B1(\mem[150][5] ), .B2(n7337), 
        .Z(n2258) );
  OA22D0 U5706 ( .A1(n7338), .A2(prog_data[4]), .B1(\mem[150][4] ), .B2(n7337), 
        .Z(n2257) );
  OA22D0 U5707 ( .A1(n7338), .A2(prog_data[3]), .B1(\mem[150][3] ), .B2(n7337), 
        .Z(n2256) );
  OA22D0 U5708 ( .A1(n7338), .A2(prog_data[2]), .B1(\mem[150][2] ), .B2(n7337), 
        .Z(n2255) );
  OA22D0 U5709 ( .A1(n7338), .A2(prog_data[1]), .B1(\mem[150][1] ), .B2(n7337), 
        .Z(n2254) );
  OA22D0 U5710 ( .A1(n7338), .A2(prog_data[0]), .B1(\mem[150][0] ), .B2(n7337), 
        .Z(n2253) );
  INVD0 U5711 ( .I(n7339), .ZN(n7340) );
  OA22D0 U5712 ( .A1(n7340), .A2(prog_data[15]), .B1(\mem[151][15] ), .B2(
        n7339), .Z(n2252) );
  OA22D0 U5713 ( .A1(n7340), .A2(prog_data[14]), .B1(\mem[151][14] ), .B2(
        n7339), .Z(n2251) );
  OA22D0 U5714 ( .A1(n7340), .A2(prog_data[13]), .B1(\mem[151][13] ), .B2(
        n7339), .Z(n2250) );
  OA22D0 U5715 ( .A1(n7340), .A2(prog_data[12]), .B1(\mem[151][12] ), .B2(
        n7339), .Z(n2249) );
  OA22D0 U5716 ( .A1(n7340), .A2(prog_data[11]), .B1(\mem[151][11] ), .B2(
        n7339), .Z(n2248) );
  OA22D0 U5717 ( .A1(n7340), .A2(prog_data[10]), .B1(\mem[151][10] ), .B2(
        n7339), .Z(n2247) );
  OA22D0 U5718 ( .A1(n7340), .A2(prog_data[9]), .B1(\mem[151][9] ), .B2(n7339), 
        .Z(n2246) );
  OA22D0 U5719 ( .A1(n7340), .A2(prog_data[8]), .B1(\mem[151][8] ), .B2(n7339), 
        .Z(n2245) );
  OA22D0 U5720 ( .A1(n7340), .A2(prog_data[7]), .B1(\mem[151][7] ), .B2(n7339), 
        .Z(n2244) );
  OA22D0 U5721 ( .A1(n7340), .A2(prog_data[6]), .B1(\mem[151][6] ), .B2(n7339), 
        .Z(n2243) );
  OA22D0 U5722 ( .A1(n7340), .A2(prog_data[5]), .B1(\mem[151][5] ), .B2(n7339), 
        .Z(n2242) );
  OA22D0 U5723 ( .A1(n7340), .A2(prog_data[4]), .B1(\mem[151][4] ), .B2(n7339), 
        .Z(n2241) );
  OA22D0 U5724 ( .A1(n7340), .A2(prog_data[3]), .B1(\mem[151][3] ), .B2(n7339), 
        .Z(n2240) );
  OA22D0 U5725 ( .A1(n7340), .A2(prog_data[2]), .B1(\mem[151][2] ), .B2(n7339), 
        .Z(n2239) );
  OA22D0 U5726 ( .A1(n7340), .A2(prog_data[1]), .B1(\mem[151][1] ), .B2(n7339), 
        .Z(n2238) );
  OA22D0 U5727 ( .A1(n7340), .A2(prog_data[0]), .B1(\mem[151][0] ), .B2(n7339), 
        .Z(n2237) );
  NR2D0 U5728 ( .A1(n7552), .A2(n7355), .ZN(n7341) );
  INVD0 U5729 ( .I(n7341), .ZN(n7342) );
  OA22D0 U5730 ( .A1(n7342), .A2(prog_data[15]), .B1(\mem[152][15] ), .B2(
        n7341), .Z(n2236) );
  OA22D0 U5731 ( .A1(n7342), .A2(prog_data[14]), .B1(\mem[152][14] ), .B2(
        n7341), .Z(n2235) );
  OA22D0 U5732 ( .A1(n7342), .A2(prog_data[13]), .B1(\mem[152][13] ), .B2(
        n7341), .Z(n2234) );
  OA22D0 U5733 ( .A1(n7342), .A2(prog_data[12]), .B1(\mem[152][12] ), .B2(
        n7341), .Z(n2233) );
  OA22D0 U5734 ( .A1(n7342), .A2(prog_data[11]), .B1(\mem[152][11] ), .B2(
        n7341), .Z(n2232) );
  OA22D0 U5735 ( .A1(n7342), .A2(prog_data[10]), .B1(\mem[152][10] ), .B2(
        n7341), .Z(n2231) );
  OA22D0 U5736 ( .A1(n7342), .A2(prog_data[9]), .B1(\mem[152][9] ), .B2(n7341), 
        .Z(n2230) );
  OA22D0 U5737 ( .A1(n7342), .A2(prog_data[8]), .B1(\mem[152][8] ), .B2(n7341), 
        .Z(n2229) );
  OA22D0 U5738 ( .A1(n7342), .A2(prog_data[7]), .B1(\mem[152][7] ), .B2(n7341), 
        .Z(n2228) );
  OA22D0 U5739 ( .A1(n7342), .A2(prog_data[6]), .B1(\mem[152][6] ), .B2(n7341), 
        .Z(n2227) );
  OA22D0 U5740 ( .A1(n7342), .A2(prog_data[5]), .B1(\mem[152][5] ), .B2(n7341), 
        .Z(n2226) );
  OA22D0 U5741 ( .A1(n7342), .A2(prog_data[4]), .B1(\mem[152][4] ), .B2(n7341), 
        .Z(n2225) );
  OA22D0 U5742 ( .A1(n7342), .A2(prog_data[3]), .B1(\mem[152][3] ), .B2(n7341), 
        .Z(n2224) );
  OA22D0 U5743 ( .A1(n7342), .A2(prog_data[2]), .B1(\mem[152][2] ), .B2(n7341), 
        .Z(n2223) );
  OA22D0 U5744 ( .A1(n7342), .A2(prog_data[1]), .B1(\mem[152][1] ), .B2(n7341), 
        .Z(n2222) );
  OA22D0 U5745 ( .A1(n7342), .A2(prog_data[0]), .B1(\mem[152][0] ), .B2(n7341), 
        .Z(n2221) );
  NR2D0 U5746 ( .A1(n7555), .A2(n7355), .ZN(n7343) );
  INVD0 U5747 ( .I(n7343), .ZN(n7344) );
  OA22D0 U5748 ( .A1(n7344), .A2(prog_data[15]), .B1(\mem[153][15] ), .B2(
        n7343), .Z(n2220) );
  OA22D0 U5749 ( .A1(n7344), .A2(prog_data[14]), .B1(\mem[153][14] ), .B2(
        n7343), .Z(n2219) );
  OA22D0 U5750 ( .A1(n7344), .A2(prog_data[13]), .B1(\mem[153][13] ), .B2(
        n7343), .Z(n2218) );
  OA22D0 U5751 ( .A1(n7344), .A2(prog_data[12]), .B1(\mem[153][12] ), .B2(
        n7343), .Z(n2217) );
  OA22D0 U5752 ( .A1(n7344), .A2(prog_data[11]), .B1(\mem[153][11] ), .B2(
        n7343), .Z(n2216) );
  OA22D0 U5753 ( .A1(n7344), .A2(prog_data[10]), .B1(\mem[153][10] ), .B2(
        n7343), .Z(n2215) );
  OA22D0 U5754 ( .A1(n7344), .A2(prog_data[9]), .B1(\mem[153][9] ), .B2(n7343), 
        .Z(n2214) );
  OA22D0 U5755 ( .A1(n7344), .A2(prog_data[8]), .B1(\mem[153][8] ), .B2(n7343), 
        .Z(n2213) );
  OA22D0 U5756 ( .A1(n7344), .A2(prog_data[7]), .B1(\mem[153][7] ), .B2(n7343), 
        .Z(n2212) );
  OA22D0 U5757 ( .A1(n7344), .A2(prog_data[6]), .B1(\mem[153][6] ), .B2(n7343), 
        .Z(n2211) );
  OA22D0 U5758 ( .A1(n7344), .A2(prog_data[5]), .B1(\mem[153][5] ), .B2(n7343), 
        .Z(n2210) );
  OA22D0 U5759 ( .A1(n7344), .A2(prog_data[4]), .B1(\mem[153][4] ), .B2(n7343), 
        .Z(n2209) );
  OA22D0 U5760 ( .A1(n7344), .A2(prog_data[3]), .B1(\mem[153][3] ), .B2(n7343), 
        .Z(n2208) );
  OA22D0 U5761 ( .A1(n7344), .A2(prog_data[2]), .B1(\mem[153][2] ), .B2(n7343), 
        .Z(n2207) );
  OA22D0 U5762 ( .A1(n7344), .A2(prog_data[1]), .B1(\mem[153][1] ), .B2(n7343), 
        .Z(n2206) );
  OA22D0 U5763 ( .A1(n7344), .A2(prog_data[0]), .B1(\mem[153][0] ), .B2(n7343), 
        .Z(n2205) );
  NR2D0 U5764 ( .A1(n7558), .A2(n7355), .ZN(n7345) );
  INVD0 U5765 ( .I(n7345), .ZN(n7346) );
  OA22D0 U5766 ( .A1(n7346), .A2(prog_data[15]), .B1(\mem[154][15] ), .B2(
        n7345), .Z(n2204) );
  OA22D0 U5767 ( .A1(n7346), .A2(prog_data[14]), .B1(\mem[154][14] ), .B2(
        n7345), .Z(n2203) );
  OA22D0 U5768 ( .A1(n7346), .A2(prog_data[13]), .B1(\mem[154][13] ), .B2(
        n7345), .Z(n2202) );
  OA22D0 U5769 ( .A1(n7346), .A2(prog_data[12]), .B1(\mem[154][12] ), .B2(
        n7345), .Z(n2201) );
  OA22D0 U5770 ( .A1(n7346), .A2(prog_data[11]), .B1(\mem[154][11] ), .B2(
        n7345), .Z(n2200) );
  OA22D0 U5771 ( .A1(n7346), .A2(prog_data[10]), .B1(\mem[154][10] ), .B2(
        n7345), .Z(n2199) );
  OA22D0 U5772 ( .A1(n7346), .A2(prog_data[9]), .B1(\mem[154][9] ), .B2(n7345), 
        .Z(n2198) );
  OA22D0 U5773 ( .A1(n7346), .A2(prog_data[8]), .B1(\mem[154][8] ), .B2(n7345), 
        .Z(n2197) );
  OA22D0 U5774 ( .A1(n7346), .A2(prog_data[7]), .B1(\mem[154][7] ), .B2(n7345), 
        .Z(n2196) );
  OA22D0 U5775 ( .A1(n7346), .A2(prog_data[6]), .B1(\mem[154][6] ), .B2(n7345), 
        .Z(n2195) );
  OA22D0 U5776 ( .A1(n7346), .A2(prog_data[5]), .B1(\mem[154][5] ), .B2(n7345), 
        .Z(n2194) );
  OA22D0 U5777 ( .A1(n7346), .A2(prog_data[4]), .B1(\mem[154][4] ), .B2(n7345), 
        .Z(n2193) );
  OA22D0 U5778 ( .A1(n7346), .A2(prog_data[3]), .B1(\mem[154][3] ), .B2(n7345), 
        .Z(n2192) );
  OA22D0 U5779 ( .A1(n7346), .A2(prog_data[2]), .B1(\mem[154][2] ), .B2(n7345), 
        .Z(n2191) );
  OA22D0 U5780 ( .A1(n7346), .A2(prog_data[1]), .B1(\mem[154][1] ), .B2(n7345), 
        .Z(n2190) );
  OA22D0 U5781 ( .A1(n7346), .A2(prog_data[0]), .B1(\mem[154][0] ), .B2(n7345), 
        .Z(n2189) );
  NR2D0 U5782 ( .A1(n7561), .A2(n7355), .ZN(n7347) );
  INVD0 U5783 ( .I(n7347), .ZN(n7348) );
  OA22D0 U5784 ( .A1(n7348), .A2(prog_data[15]), .B1(\mem[155][15] ), .B2(
        n7347), .Z(n2188) );
  OA22D0 U5785 ( .A1(n7348), .A2(prog_data[14]), .B1(\mem[155][14] ), .B2(
        n7347), .Z(n2187) );
  OA22D0 U5786 ( .A1(n7348), .A2(prog_data[13]), .B1(\mem[155][13] ), .B2(
        n7347), .Z(n2186) );
  OA22D0 U5787 ( .A1(n7348), .A2(prog_data[12]), .B1(\mem[155][12] ), .B2(
        n7347), .Z(n2185) );
  OA22D0 U5788 ( .A1(n7348), .A2(prog_data[11]), .B1(\mem[155][11] ), .B2(
        n7347), .Z(n2184) );
  OA22D0 U5789 ( .A1(n7348), .A2(prog_data[10]), .B1(\mem[155][10] ), .B2(
        n7347), .Z(n2183) );
  OA22D0 U5790 ( .A1(n7348), .A2(prog_data[9]), .B1(\mem[155][9] ), .B2(n7347), 
        .Z(n2182) );
  OA22D0 U5791 ( .A1(n7348), .A2(prog_data[8]), .B1(\mem[155][8] ), .B2(n7347), 
        .Z(n2181) );
  OA22D0 U5792 ( .A1(n7348), .A2(prog_data[7]), .B1(\mem[155][7] ), .B2(n7347), 
        .Z(n2180) );
  OA22D0 U5793 ( .A1(n7348), .A2(prog_data[6]), .B1(\mem[155][6] ), .B2(n7347), 
        .Z(n2179) );
  OA22D0 U5794 ( .A1(n7348), .A2(prog_data[5]), .B1(\mem[155][5] ), .B2(n7347), 
        .Z(n2178) );
  OA22D0 U5795 ( .A1(n7348), .A2(prog_data[4]), .B1(\mem[155][4] ), .B2(n7347), 
        .Z(n2177) );
  OA22D0 U5796 ( .A1(n7348), .A2(prog_data[3]), .B1(\mem[155][3] ), .B2(n7347), 
        .Z(n2176) );
  OA22D0 U5797 ( .A1(n7348), .A2(prog_data[2]), .B1(\mem[155][2] ), .B2(n7347), 
        .Z(n2175) );
  OA22D0 U5798 ( .A1(n7348), .A2(prog_data[1]), .B1(\mem[155][1] ), .B2(n7347), 
        .Z(n2174) );
  OA22D0 U5799 ( .A1(n7348), .A2(prog_data[0]), .B1(\mem[155][0] ), .B2(n7347), 
        .Z(n2173) );
  NR2D0 U5800 ( .A1(n7564), .A2(n7355), .ZN(n7349) );
  INVD0 U5801 ( .I(n7349), .ZN(n7350) );
  OA22D0 U5802 ( .A1(n7350), .A2(prog_data[15]), .B1(\mem[156][15] ), .B2(
        n7349), .Z(n2172) );
  OA22D0 U5803 ( .A1(n7350), .A2(prog_data[14]), .B1(\mem[156][14] ), .B2(
        n7349), .Z(n2171) );
  OA22D0 U5804 ( .A1(n7350), .A2(prog_data[13]), .B1(\mem[156][13] ), .B2(
        n7349), .Z(n2170) );
  OA22D0 U5805 ( .A1(n7350), .A2(prog_data[12]), .B1(\mem[156][12] ), .B2(
        n7349), .Z(n2169) );
  OA22D0 U5806 ( .A1(n7350), .A2(prog_data[11]), .B1(\mem[156][11] ), .B2(
        n7349), .Z(n2168) );
  OA22D0 U5807 ( .A1(n7350), .A2(prog_data[10]), .B1(\mem[156][10] ), .B2(
        n7349), .Z(n2167) );
  OA22D0 U5808 ( .A1(n7350), .A2(prog_data[9]), .B1(\mem[156][9] ), .B2(n7349), 
        .Z(n2166) );
  OA22D0 U5809 ( .A1(n7350), .A2(prog_data[8]), .B1(\mem[156][8] ), .B2(n7349), 
        .Z(n2165) );
  OA22D0 U5810 ( .A1(n7350), .A2(prog_data[7]), .B1(\mem[156][7] ), .B2(n7349), 
        .Z(n2164) );
  OA22D0 U5811 ( .A1(n7350), .A2(prog_data[6]), .B1(\mem[156][6] ), .B2(n7349), 
        .Z(n2163) );
  OA22D0 U5812 ( .A1(n7350), .A2(prog_data[5]), .B1(\mem[156][5] ), .B2(n7349), 
        .Z(n2162) );
  OA22D0 U5813 ( .A1(n7350), .A2(prog_data[4]), .B1(\mem[156][4] ), .B2(n7349), 
        .Z(n2161) );
  OA22D0 U5814 ( .A1(n7350), .A2(prog_data[3]), .B1(\mem[156][3] ), .B2(n7349), 
        .Z(n2160) );
  OA22D0 U5815 ( .A1(n7350), .A2(prog_data[2]), .B1(\mem[156][2] ), .B2(n7349), 
        .Z(n2159) );
  OA22D0 U5816 ( .A1(n7350), .A2(prog_data[1]), .B1(\mem[156][1] ), .B2(n7349), 
        .Z(n2158) );
  OA22D0 U5817 ( .A1(n7350), .A2(prog_data[0]), .B1(\mem[156][0] ), .B2(n7349), 
        .Z(n2157) );
  NR2D0 U5818 ( .A1(n7567), .A2(n7355), .ZN(n7351) );
  INVD0 U5819 ( .I(n7351), .ZN(n7352) );
  OA22D0 U5820 ( .A1(n7352), .A2(prog_data[15]), .B1(\mem[157][15] ), .B2(
        n7351), .Z(n2156) );
  OA22D0 U5821 ( .A1(n7352), .A2(prog_data[14]), .B1(\mem[157][14] ), .B2(
        n7351), .Z(n2155) );
  OA22D0 U5822 ( .A1(n7352), .A2(prog_data[13]), .B1(\mem[157][13] ), .B2(
        n7351), .Z(n2154) );
  OA22D0 U5823 ( .A1(n7352), .A2(prog_data[12]), .B1(\mem[157][12] ), .B2(
        n7351), .Z(n2153) );
  OA22D0 U5824 ( .A1(n7352), .A2(prog_data[11]), .B1(\mem[157][11] ), .B2(
        n7351), .Z(n2152) );
  OA22D0 U5825 ( .A1(n7352), .A2(prog_data[10]), .B1(\mem[157][10] ), .B2(
        n7351), .Z(n2151) );
  OA22D0 U5826 ( .A1(n7352), .A2(prog_data[9]), .B1(\mem[157][9] ), .B2(n7351), 
        .Z(n2150) );
  OA22D0 U5827 ( .A1(n7352), .A2(prog_data[8]), .B1(\mem[157][8] ), .B2(n7351), 
        .Z(n2149) );
  OA22D0 U5828 ( .A1(n7352), .A2(prog_data[7]), .B1(\mem[157][7] ), .B2(n7351), 
        .Z(n2148) );
  OA22D0 U5829 ( .A1(n7352), .A2(prog_data[6]), .B1(\mem[157][6] ), .B2(n7351), 
        .Z(n2147) );
  OA22D0 U5830 ( .A1(n7352), .A2(prog_data[5]), .B1(\mem[157][5] ), .B2(n7351), 
        .Z(n2146) );
  OA22D0 U5831 ( .A1(n7352), .A2(prog_data[4]), .B1(\mem[157][4] ), .B2(n7351), 
        .Z(n2145) );
  OA22D0 U5832 ( .A1(n7352), .A2(prog_data[3]), .B1(\mem[157][3] ), .B2(n7351), 
        .Z(n2144) );
  OA22D0 U5833 ( .A1(n7352), .A2(prog_data[2]), .B1(\mem[157][2] ), .B2(n7351), 
        .Z(n2143) );
  OA22D0 U5834 ( .A1(n7352), .A2(prog_data[1]), .B1(\mem[157][1] ), .B2(n7351), 
        .Z(n2142) );
  OA22D0 U5835 ( .A1(n7352), .A2(prog_data[0]), .B1(\mem[157][0] ), .B2(n7351), 
        .Z(n2141) );
  NR2D0 U5836 ( .A1(n7570), .A2(n7355), .ZN(n7353) );
  INVD0 U5837 ( .I(n7353), .ZN(n7354) );
  OA22D0 U5838 ( .A1(n7354), .A2(prog_data[15]), .B1(\mem[158][15] ), .B2(
        n7353), .Z(n2140) );
  OA22D0 U5839 ( .A1(n7354), .A2(prog_data[14]), .B1(\mem[158][14] ), .B2(
        n7353), .Z(n2139) );
  OA22D0 U5840 ( .A1(n7354), .A2(prog_data[13]), .B1(\mem[158][13] ), .B2(
        n7353), .Z(n2138) );
  OA22D0 U5841 ( .A1(n7354), .A2(prog_data[12]), .B1(\mem[158][12] ), .B2(
        n7353), .Z(n2137) );
  OA22D0 U5842 ( .A1(n7354), .A2(prog_data[11]), .B1(\mem[158][11] ), .B2(
        n7353), .Z(n2136) );
  OA22D0 U5843 ( .A1(n7354), .A2(prog_data[10]), .B1(\mem[158][10] ), .B2(
        n7353), .Z(n2135) );
  OA22D0 U5844 ( .A1(n7354), .A2(prog_data[9]), .B1(\mem[158][9] ), .B2(n7353), 
        .Z(n2134) );
  OA22D0 U5845 ( .A1(n7354), .A2(prog_data[8]), .B1(\mem[158][8] ), .B2(n7353), 
        .Z(n2133) );
  OA22D0 U5846 ( .A1(n7354), .A2(prog_data[7]), .B1(\mem[158][7] ), .B2(n7353), 
        .Z(n2132) );
  OA22D0 U5847 ( .A1(n7354), .A2(prog_data[6]), .B1(\mem[158][6] ), .B2(n7353), 
        .Z(n2131) );
  OA22D0 U5848 ( .A1(n7354), .A2(prog_data[5]), .B1(\mem[158][5] ), .B2(n7353), 
        .Z(n2130) );
  OA22D0 U5849 ( .A1(n7354), .A2(prog_data[4]), .B1(\mem[158][4] ), .B2(n7353), 
        .Z(n2129) );
  OA22D0 U5850 ( .A1(n7354), .A2(prog_data[3]), .B1(\mem[158][3] ), .B2(n7353), 
        .Z(n2128) );
  OA22D0 U5851 ( .A1(n7354), .A2(prog_data[2]), .B1(\mem[158][2] ), .B2(n7353), 
        .Z(n2127) );
  OA22D0 U5852 ( .A1(n7354), .A2(prog_data[1]), .B1(\mem[158][1] ), .B2(n7353), 
        .Z(n2126) );
  OA22D0 U5853 ( .A1(n7354), .A2(prog_data[0]), .B1(\mem[158][0] ), .B2(n7353), 
        .Z(n2125) );
  NR2D0 U5854 ( .A1(n7574), .A2(n7355), .ZN(n7356) );
  OA22D0 U5855 ( .A1(n7357), .A2(prog_data[15]), .B1(\mem[159][15] ), .B2(
        n7356), .Z(n2124) );
  OA22D0 U5856 ( .A1(n7357), .A2(prog_data[14]), .B1(\mem[159][14] ), .B2(
        n7356), .Z(n2123) );
  OA22D0 U5857 ( .A1(n7357), .A2(prog_data[13]), .B1(\mem[159][13] ), .B2(
        n7356), .Z(n2122) );
  OA22D0 U5858 ( .A1(n7357), .A2(prog_data[12]), .B1(\mem[159][12] ), .B2(
        n7356), .Z(n2121) );
  OA22D0 U5859 ( .A1(n7357), .A2(prog_data[11]), .B1(\mem[159][11] ), .B2(
        n7356), .Z(n2120) );
  OA22D0 U5860 ( .A1(n7357), .A2(prog_data[10]), .B1(\mem[159][10] ), .B2(
        n7356), .Z(n2119) );
  OA22D0 U5861 ( .A1(n7357), .A2(prog_data[9]), .B1(\mem[159][9] ), .B2(n7356), 
        .Z(n2118) );
  OA22D0 U5862 ( .A1(n7357), .A2(prog_data[8]), .B1(\mem[159][8] ), .B2(n7356), 
        .Z(n2117) );
  OA22D0 U5863 ( .A1(n7357), .A2(prog_data[7]), .B1(\mem[159][7] ), .B2(n7356), 
        .Z(n2116) );
  OA22D0 U5864 ( .A1(n7357), .A2(prog_data[6]), .B1(\mem[159][6] ), .B2(n7356), 
        .Z(n2115) );
  OA22D0 U5865 ( .A1(n7357), .A2(prog_data[5]), .B1(\mem[159][5] ), .B2(n7356), 
        .Z(n2114) );
  OA22D0 U5866 ( .A1(n7357), .A2(prog_data[4]), .B1(\mem[159][4] ), .B2(n7356), 
        .Z(n2113) );
  OA22D0 U5867 ( .A1(n7357), .A2(prog_data[3]), .B1(\mem[159][3] ), .B2(n7356), 
        .Z(n2112) );
  OA22D0 U5868 ( .A1(n7357), .A2(prog_data[2]), .B1(\mem[159][2] ), .B2(n7356), 
        .Z(n2111) );
  OA22D0 U5869 ( .A1(n7357), .A2(prog_data[1]), .B1(\mem[159][1] ), .B2(n7356), 
        .Z(n2110) );
  OA22D0 U5870 ( .A1(n7357), .A2(prog_data[0]), .B1(\mem[159][0] ), .B2(n7356), 
        .Z(n2109) );
  CKND2D0 U5871 ( .A1(prog_addr[5]), .A2(prog_we), .ZN(n7527) );
  CKND2D0 U5872 ( .A1(n7492), .A2(n7391), .ZN(n7388) );
  NR2D0 U5873 ( .A1(n7528), .A2(n7388), .ZN(n7358) );
  INVD0 U5874 ( .I(n7358), .ZN(n7359) );
  OA22D0 U5875 ( .A1(n7359), .A2(prog_data[15]), .B1(\mem[160][15] ), .B2(
        n7358), .Z(n2108) );
  OA22D0 U5876 ( .A1(n7359), .A2(prog_data[14]), .B1(\mem[160][14] ), .B2(
        n7358), .Z(n2107) );
  OA22D0 U5877 ( .A1(n7359), .A2(prog_data[13]), .B1(\mem[160][13] ), .B2(
        n7358), .Z(n2106) );
  OA22D0 U5878 ( .A1(n7359), .A2(prog_data[12]), .B1(\mem[160][12] ), .B2(
        n7358), .Z(n2105) );
  OA22D0 U5879 ( .A1(n7359), .A2(prog_data[11]), .B1(\mem[160][11] ), .B2(
        n7358), .Z(n2104) );
  OA22D0 U5880 ( .A1(n7359), .A2(prog_data[10]), .B1(\mem[160][10] ), .B2(
        n7358), .Z(n2103) );
  OA22D0 U5881 ( .A1(n7359), .A2(prog_data[9]), .B1(\mem[160][9] ), .B2(n7358), 
        .Z(n2102) );
  OA22D0 U5882 ( .A1(n7359), .A2(prog_data[8]), .B1(\mem[160][8] ), .B2(n7358), 
        .Z(n2101) );
  OA22D0 U5883 ( .A1(n7359), .A2(prog_data[7]), .B1(\mem[160][7] ), .B2(n7358), 
        .Z(n2100) );
  OA22D0 U5884 ( .A1(n7359), .A2(prog_data[6]), .B1(\mem[160][6] ), .B2(n7358), 
        .Z(n2099) );
  OA22D0 U5885 ( .A1(n7359), .A2(prog_data[5]), .B1(\mem[160][5] ), .B2(n7358), 
        .Z(n2098) );
  OA22D0 U5886 ( .A1(n7359), .A2(prog_data[4]), .B1(\mem[160][4] ), .B2(n7358), 
        .Z(n2097) );
  OA22D0 U5887 ( .A1(n7359), .A2(prog_data[3]), .B1(\mem[160][3] ), .B2(n7358), 
        .Z(n2096) );
  OA22D0 U5888 ( .A1(n7359), .A2(prog_data[2]), .B1(\mem[160][2] ), .B2(n7358), 
        .Z(n2095) );
  OA22D0 U5889 ( .A1(n7359), .A2(prog_data[1]), .B1(\mem[160][1] ), .B2(n7358), 
        .Z(n2094) );
  OA22D0 U5890 ( .A1(n7359), .A2(prog_data[0]), .B1(\mem[160][0] ), .B2(n7358), 
        .Z(n2093) );
  NR2D0 U5891 ( .A1(n7531), .A2(n7388), .ZN(n7360) );
  INVD0 U5892 ( .I(n7360), .ZN(n7361) );
  OA22D0 U5893 ( .A1(n7361), .A2(prog_data[15]), .B1(\mem[161][15] ), .B2(
        n7360), .Z(n2092) );
  OA22D0 U5894 ( .A1(n7361), .A2(prog_data[14]), .B1(\mem[161][14] ), .B2(
        n7360), .Z(n2091) );
  OA22D0 U5895 ( .A1(n7361), .A2(prog_data[13]), .B1(\mem[161][13] ), .B2(
        n7360), .Z(n2090) );
  OA22D0 U5896 ( .A1(n7361), .A2(prog_data[12]), .B1(\mem[161][12] ), .B2(
        n7360), .Z(n2089) );
  OA22D0 U5897 ( .A1(n7361), .A2(prog_data[11]), .B1(\mem[161][11] ), .B2(
        n7360), .Z(n2088) );
  OA22D0 U5898 ( .A1(n7361), .A2(prog_data[10]), .B1(\mem[161][10] ), .B2(
        n7360), .Z(n2087) );
  OA22D0 U5899 ( .A1(n7361), .A2(prog_data[9]), .B1(\mem[161][9] ), .B2(n7360), 
        .Z(n2086) );
  OA22D0 U5900 ( .A1(n7361), .A2(prog_data[8]), .B1(\mem[161][8] ), .B2(n7360), 
        .Z(n2085) );
  OA22D0 U5901 ( .A1(n7361), .A2(prog_data[7]), .B1(\mem[161][7] ), .B2(n7360), 
        .Z(n2084) );
  OA22D0 U5902 ( .A1(n7361), .A2(prog_data[6]), .B1(\mem[161][6] ), .B2(n7360), 
        .Z(n2083) );
  OA22D0 U5903 ( .A1(n7361), .A2(prog_data[5]), .B1(\mem[161][5] ), .B2(n7360), 
        .Z(n2082) );
  OA22D0 U5904 ( .A1(n7361), .A2(prog_data[4]), .B1(\mem[161][4] ), .B2(n7360), 
        .Z(n2081) );
  OA22D0 U5905 ( .A1(n7361), .A2(prog_data[3]), .B1(\mem[161][3] ), .B2(n7360), 
        .Z(n2080) );
  OA22D0 U5906 ( .A1(n7361), .A2(prog_data[2]), .B1(\mem[161][2] ), .B2(n7360), 
        .Z(n2079) );
  OA22D0 U5907 ( .A1(n7361), .A2(prog_data[1]), .B1(\mem[161][1] ), .B2(n7360), 
        .Z(n2078) );
  OA22D0 U5908 ( .A1(n7361), .A2(prog_data[0]), .B1(\mem[161][0] ), .B2(n7360), 
        .Z(n2077) );
  NR2D0 U5909 ( .A1(n7534), .A2(n7388), .ZN(n7362) );
  INVD0 U5910 ( .I(n7362), .ZN(n7363) );
  OA22D0 U5911 ( .A1(n7363), .A2(prog_data[15]), .B1(\mem[162][15] ), .B2(
        n7362), .Z(n2076) );
  OA22D0 U5912 ( .A1(n7363), .A2(prog_data[14]), .B1(\mem[162][14] ), .B2(
        n7362), .Z(n2075) );
  OA22D0 U5913 ( .A1(n7363), .A2(prog_data[13]), .B1(\mem[162][13] ), .B2(
        n7362), .Z(n2074) );
  OA22D0 U5914 ( .A1(n7363), .A2(prog_data[12]), .B1(\mem[162][12] ), .B2(
        n7362), .Z(n2073) );
  OA22D0 U5915 ( .A1(n7363), .A2(prog_data[11]), .B1(\mem[162][11] ), .B2(
        n7362), .Z(n2072) );
  OA22D0 U5916 ( .A1(n7363), .A2(prog_data[10]), .B1(\mem[162][10] ), .B2(
        n7362), .Z(n2071) );
  OA22D0 U5917 ( .A1(n7363), .A2(prog_data[9]), .B1(\mem[162][9] ), .B2(n7362), 
        .Z(n2070) );
  OA22D0 U5918 ( .A1(n7363), .A2(prog_data[8]), .B1(\mem[162][8] ), .B2(n7362), 
        .Z(n2069) );
  OA22D0 U5919 ( .A1(n7363), .A2(prog_data[7]), .B1(\mem[162][7] ), .B2(n7362), 
        .Z(n2068) );
  OA22D0 U5920 ( .A1(n7363), .A2(prog_data[6]), .B1(\mem[162][6] ), .B2(n7362), 
        .Z(n2067) );
  OA22D0 U5921 ( .A1(n7363), .A2(prog_data[5]), .B1(\mem[162][5] ), .B2(n7362), 
        .Z(n2066) );
  OA22D0 U5922 ( .A1(n7363), .A2(prog_data[4]), .B1(\mem[162][4] ), .B2(n7362), 
        .Z(n2065) );
  OA22D0 U5923 ( .A1(n7363), .A2(prog_data[3]), .B1(\mem[162][3] ), .B2(n7362), 
        .Z(n2064) );
  OA22D0 U5924 ( .A1(n7363), .A2(prog_data[2]), .B1(\mem[162][2] ), .B2(n7362), 
        .Z(n2063) );
  OA22D0 U5925 ( .A1(n7363), .A2(prog_data[1]), .B1(\mem[162][1] ), .B2(n7362), 
        .Z(n2062) );
  OA22D0 U5926 ( .A1(n7363), .A2(prog_data[0]), .B1(\mem[162][0] ), .B2(n7362), 
        .Z(n2061) );
  NR2D0 U5927 ( .A1(n7537), .A2(n7388), .ZN(n7364) );
  INVD0 U5928 ( .I(n7364), .ZN(n7365) );
  OA22D0 U5929 ( .A1(n7365), .A2(prog_data[15]), .B1(\mem[163][15] ), .B2(
        n7364), .Z(n2060) );
  OA22D0 U5930 ( .A1(n7365), .A2(prog_data[14]), .B1(\mem[163][14] ), .B2(
        n7364), .Z(n2059) );
  OA22D0 U5931 ( .A1(n7365), .A2(prog_data[13]), .B1(\mem[163][13] ), .B2(
        n7364), .Z(n2058) );
  OA22D0 U5932 ( .A1(n7365), .A2(prog_data[12]), .B1(\mem[163][12] ), .B2(
        n7364), .Z(n2057) );
  OA22D0 U5933 ( .A1(n7365), .A2(prog_data[11]), .B1(\mem[163][11] ), .B2(
        n7364), .Z(n2056) );
  OA22D0 U5934 ( .A1(n7365), .A2(prog_data[10]), .B1(\mem[163][10] ), .B2(
        n7364), .Z(n2055) );
  OA22D0 U5935 ( .A1(n7365), .A2(prog_data[9]), .B1(\mem[163][9] ), .B2(n7364), 
        .Z(n2054) );
  OA22D0 U5936 ( .A1(n7365), .A2(prog_data[8]), .B1(\mem[163][8] ), .B2(n7364), 
        .Z(n2053) );
  OA22D0 U5937 ( .A1(n7365), .A2(prog_data[7]), .B1(\mem[163][7] ), .B2(n7364), 
        .Z(n2052) );
  OA22D0 U5938 ( .A1(n7365), .A2(prog_data[6]), .B1(\mem[163][6] ), .B2(n7364), 
        .Z(n2051) );
  OA22D0 U5939 ( .A1(n7365), .A2(prog_data[5]), .B1(\mem[163][5] ), .B2(n7364), 
        .Z(n2050) );
  OA22D0 U5940 ( .A1(n7365), .A2(prog_data[4]), .B1(\mem[163][4] ), .B2(n7364), 
        .Z(n2049) );
  OA22D0 U5941 ( .A1(n7365), .A2(prog_data[3]), .B1(\mem[163][3] ), .B2(n7364), 
        .Z(n2048) );
  OA22D0 U5942 ( .A1(n7365), .A2(prog_data[2]), .B1(\mem[163][2] ), .B2(n7364), 
        .Z(n2047) );
  OA22D0 U5943 ( .A1(n7365), .A2(prog_data[1]), .B1(\mem[163][1] ), .B2(n7364), 
        .Z(n2046) );
  OA22D0 U5944 ( .A1(n7365), .A2(prog_data[0]), .B1(\mem[163][0] ), .B2(n7364), 
        .Z(n2045) );
  NR2D0 U5945 ( .A1(n7540), .A2(n7388), .ZN(n7366) );
  INVD0 U5946 ( .I(n7366), .ZN(n7367) );
  OA22D0 U5947 ( .A1(n7367), .A2(prog_data[15]), .B1(\mem[164][15] ), .B2(
        n7366), .Z(n2044) );
  OA22D0 U5948 ( .A1(n7367), .A2(prog_data[14]), .B1(\mem[164][14] ), .B2(
        n7366), .Z(n2043) );
  OA22D0 U5949 ( .A1(n7367), .A2(prog_data[13]), .B1(\mem[164][13] ), .B2(
        n7366), .Z(n2042) );
  OA22D0 U5950 ( .A1(n7367), .A2(prog_data[12]), .B1(\mem[164][12] ), .B2(
        n7366), .Z(n2041) );
  OA22D0 U5951 ( .A1(n7367), .A2(prog_data[11]), .B1(\mem[164][11] ), .B2(
        n7366), .Z(n2040) );
  OA22D0 U5952 ( .A1(n7367), .A2(prog_data[10]), .B1(\mem[164][10] ), .B2(
        n7366), .Z(n2039) );
  OA22D0 U5953 ( .A1(n7367), .A2(prog_data[9]), .B1(\mem[164][9] ), .B2(n7366), 
        .Z(n2038) );
  OA22D0 U5954 ( .A1(n7367), .A2(prog_data[8]), .B1(\mem[164][8] ), .B2(n7366), 
        .Z(n2037) );
  OA22D0 U5955 ( .A1(n7367), .A2(prog_data[7]), .B1(\mem[164][7] ), .B2(n7366), 
        .Z(n2036) );
  OA22D0 U5956 ( .A1(n7367), .A2(prog_data[6]), .B1(\mem[164][6] ), .B2(n7366), 
        .Z(n2035) );
  OA22D0 U5957 ( .A1(n7367), .A2(prog_data[5]), .B1(\mem[164][5] ), .B2(n7366), 
        .Z(n2034) );
  OA22D0 U5958 ( .A1(n7367), .A2(prog_data[4]), .B1(\mem[164][4] ), .B2(n7366), 
        .Z(n2033) );
  OA22D0 U5959 ( .A1(n7367), .A2(prog_data[3]), .B1(\mem[164][3] ), .B2(n7366), 
        .Z(n2032) );
  OA22D0 U5960 ( .A1(n7367), .A2(prog_data[2]), .B1(\mem[164][2] ), .B2(n7366), 
        .Z(n2031) );
  OA22D0 U5961 ( .A1(n7367), .A2(prog_data[1]), .B1(\mem[164][1] ), .B2(n7366), 
        .Z(n2030) );
  OA22D0 U5962 ( .A1(n7367), .A2(prog_data[0]), .B1(\mem[164][0] ), .B2(n7366), 
        .Z(n2029) );
  NR2D0 U5963 ( .A1(n7543), .A2(n7388), .ZN(n7368) );
  INVD0 U5964 ( .I(n7368), .ZN(n7369) );
  OA22D0 U5965 ( .A1(n7369), .A2(prog_data[15]), .B1(\mem[165][15] ), .B2(
        n7368), .Z(n2028) );
  OA22D0 U5966 ( .A1(n7369), .A2(prog_data[14]), .B1(\mem[165][14] ), .B2(
        n7368), .Z(n2027) );
  OA22D0 U5967 ( .A1(n7369), .A2(prog_data[13]), .B1(\mem[165][13] ), .B2(
        n7368), .Z(n2026) );
  OA22D0 U5968 ( .A1(n7369), .A2(prog_data[12]), .B1(\mem[165][12] ), .B2(
        n7368), .Z(n2025) );
  OA22D0 U5969 ( .A1(n7369), .A2(prog_data[11]), .B1(\mem[165][11] ), .B2(
        n7368), .Z(n2024) );
  OA22D0 U5970 ( .A1(n7369), .A2(prog_data[10]), .B1(\mem[165][10] ), .B2(
        n7368), .Z(n2023) );
  OA22D0 U5971 ( .A1(n7369), .A2(prog_data[9]), .B1(\mem[165][9] ), .B2(n7368), 
        .Z(n2022) );
  OA22D0 U5972 ( .A1(n7369), .A2(prog_data[8]), .B1(\mem[165][8] ), .B2(n7368), 
        .Z(n2021) );
  OA22D0 U5973 ( .A1(n7369), .A2(prog_data[7]), .B1(\mem[165][7] ), .B2(n7368), 
        .Z(n2020) );
  OA22D0 U5974 ( .A1(n7369), .A2(prog_data[6]), .B1(\mem[165][6] ), .B2(n7368), 
        .Z(n2019) );
  OA22D0 U5975 ( .A1(n7369), .A2(prog_data[5]), .B1(\mem[165][5] ), .B2(n7368), 
        .Z(n2018) );
  OA22D0 U5976 ( .A1(n7369), .A2(prog_data[4]), .B1(\mem[165][4] ), .B2(n7368), 
        .Z(n2017) );
  OA22D0 U5977 ( .A1(n7369), .A2(prog_data[3]), .B1(\mem[165][3] ), .B2(n7368), 
        .Z(n2016) );
  OA22D0 U5978 ( .A1(n7369), .A2(prog_data[2]), .B1(\mem[165][2] ), .B2(n7368), 
        .Z(n2015) );
  OA22D0 U5979 ( .A1(n7369), .A2(prog_data[1]), .B1(\mem[165][1] ), .B2(n7368), 
        .Z(n2014) );
  OA22D0 U5980 ( .A1(n7369), .A2(prog_data[0]), .B1(\mem[165][0] ), .B2(n7368), 
        .Z(n2013) );
  INVD0 U5981 ( .I(n7370), .ZN(n7371) );
  OA22D0 U5982 ( .A1(n7371), .A2(prog_data[15]), .B1(\mem[166][15] ), .B2(
        n7370), .Z(n2012) );
  OA22D0 U5983 ( .A1(n7371), .A2(prog_data[14]), .B1(\mem[166][14] ), .B2(
        n7370), .Z(n2011) );
  OA22D0 U5984 ( .A1(n7371), .A2(prog_data[13]), .B1(\mem[166][13] ), .B2(
        n7370), .Z(n2010) );
  OA22D0 U5985 ( .A1(n7371), .A2(prog_data[12]), .B1(\mem[166][12] ), .B2(
        n7370), .Z(n2009) );
  OA22D0 U5986 ( .A1(n7371), .A2(prog_data[11]), .B1(\mem[166][11] ), .B2(
        n7370), .Z(n2008) );
  OA22D0 U5987 ( .A1(n7371), .A2(prog_data[10]), .B1(\mem[166][10] ), .B2(
        n7370), .Z(n2007) );
  OA22D0 U5988 ( .A1(n7371), .A2(prog_data[9]), .B1(\mem[166][9] ), .B2(n7370), 
        .Z(n2006) );
  OA22D0 U5989 ( .A1(n7371), .A2(prog_data[8]), .B1(\mem[166][8] ), .B2(n7370), 
        .Z(n2005) );
  OA22D0 U5990 ( .A1(n7371), .A2(prog_data[7]), .B1(\mem[166][7] ), .B2(n7370), 
        .Z(n2004) );
  OA22D0 U5991 ( .A1(n7371), .A2(prog_data[6]), .B1(\mem[166][6] ), .B2(n7370), 
        .Z(n2003) );
  OA22D0 U5992 ( .A1(n7371), .A2(prog_data[5]), .B1(\mem[166][5] ), .B2(n7370), 
        .Z(n2002) );
  OA22D0 U5993 ( .A1(n7371), .A2(prog_data[4]), .B1(\mem[166][4] ), .B2(n7370), 
        .Z(n2001) );
  OA22D0 U5994 ( .A1(n7371), .A2(prog_data[3]), .B1(\mem[166][3] ), .B2(n7370), 
        .Z(n2000) );
  OA22D0 U5995 ( .A1(n7371), .A2(prog_data[2]), .B1(\mem[166][2] ), .B2(n7370), 
        .Z(n1999) );
  OA22D0 U5996 ( .A1(n7371), .A2(prog_data[1]), .B1(\mem[166][1] ), .B2(n7370), 
        .Z(n1998) );
  OA22D0 U5997 ( .A1(n7371), .A2(prog_data[0]), .B1(\mem[166][0] ), .B2(n7370), 
        .Z(n1997) );
  NR2D0 U5998 ( .A1(n7549), .A2(n7388), .ZN(n7372) );
  INVD0 U5999 ( .I(n7372), .ZN(n7373) );
  OA22D0 U6000 ( .A1(n7373), .A2(prog_data[15]), .B1(\mem[167][15] ), .B2(
        n7372), .Z(n1996) );
  OA22D0 U6001 ( .A1(n7373), .A2(prog_data[14]), .B1(\mem[167][14] ), .B2(
        n7372), .Z(n1995) );
  OA22D0 U6002 ( .A1(n7373), .A2(prog_data[13]), .B1(\mem[167][13] ), .B2(
        n7372), .Z(n1994) );
  OA22D0 U6003 ( .A1(n7373), .A2(prog_data[12]), .B1(\mem[167][12] ), .B2(
        n7372), .Z(n1993) );
  OA22D0 U6004 ( .A1(n7373), .A2(prog_data[11]), .B1(\mem[167][11] ), .B2(
        n7372), .Z(n1992) );
  OA22D0 U6005 ( .A1(n7373), .A2(prog_data[10]), .B1(\mem[167][10] ), .B2(
        n7372), .Z(n1991) );
  OA22D0 U6006 ( .A1(n7373), .A2(prog_data[9]), .B1(\mem[167][9] ), .B2(n7372), 
        .Z(n1990) );
  OA22D0 U6007 ( .A1(n7373), .A2(prog_data[8]), .B1(\mem[167][8] ), .B2(n7372), 
        .Z(n1989) );
  OA22D0 U6008 ( .A1(n7373), .A2(prog_data[7]), .B1(\mem[167][7] ), .B2(n7372), 
        .Z(n1988) );
  OA22D0 U6009 ( .A1(n7373), .A2(prog_data[6]), .B1(\mem[167][6] ), .B2(n7372), 
        .Z(n1987) );
  OA22D0 U6010 ( .A1(n7373), .A2(prog_data[5]), .B1(\mem[167][5] ), .B2(n7372), 
        .Z(n1986) );
  OA22D0 U6011 ( .A1(n7373), .A2(prog_data[4]), .B1(\mem[167][4] ), .B2(n7372), 
        .Z(n1985) );
  OA22D0 U6012 ( .A1(n7373), .A2(prog_data[3]), .B1(\mem[167][3] ), .B2(n7372), 
        .Z(n1984) );
  OA22D0 U6013 ( .A1(n7373), .A2(prog_data[2]), .B1(\mem[167][2] ), .B2(n7372), 
        .Z(n1983) );
  OA22D0 U6014 ( .A1(n7373), .A2(prog_data[1]), .B1(\mem[167][1] ), .B2(n7372), 
        .Z(n1982) );
  OA22D0 U6015 ( .A1(n7373), .A2(prog_data[0]), .B1(\mem[167][0] ), .B2(n7372), 
        .Z(n1981) );
  NR2D0 U6016 ( .A1(n7552), .A2(n7388), .ZN(n7374) );
  INVD0 U6017 ( .I(n7374), .ZN(n7375) );
  OA22D0 U6018 ( .A1(n7375), .A2(prog_data[15]), .B1(\mem[168][15] ), .B2(
        n7374), .Z(n1980) );
  OA22D0 U6019 ( .A1(n7375), .A2(prog_data[14]), .B1(\mem[168][14] ), .B2(
        n7374), .Z(n1979) );
  OA22D0 U6020 ( .A1(n7375), .A2(prog_data[13]), .B1(\mem[168][13] ), .B2(
        n7374), .Z(n1978) );
  OA22D0 U6021 ( .A1(n7375), .A2(prog_data[12]), .B1(\mem[168][12] ), .B2(
        n7374), .Z(n1977) );
  OA22D0 U6022 ( .A1(n7375), .A2(prog_data[11]), .B1(\mem[168][11] ), .B2(
        n7374), .Z(n1976) );
  OA22D0 U6023 ( .A1(n7375), .A2(prog_data[10]), .B1(\mem[168][10] ), .B2(
        n7374), .Z(n1975) );
  OA22D0 U6024 ( .A1(n7375), .A2(prog_data[9]), .B1(\mem[168][9] ), .B2(n7374), 
        .Z(n1974) );
  OA22D0 U6025 ( .A1(n7375), .A2(prog_data[8]), .B1(\mem[168][8] ), .B2(n7374), 
        .Z(n1973) );
  OA22D0 U6026 ( .A1(n7375), .A2(prog_data[7]), .B1(\mem[168][7] ), .B2(n7374), 
        .Z(n1972) );
  OA22D0 U6027 ( .A1(n7375), .A2(prog_data[6]), .B1(\mem[168][6] ), .B2(n7374), 
        .Z(n1971) );
  OA22D0 U6028 ( .A1(n7375), .A2(prog_data[5]), .B1(\mem[168][5] ), .B2(n7374), 
        .Z(n1970) );
  OA22D0 U6029 ( .A1(n7375), .A2(prog_data[4]), .B1(\mem[168][4] ), .B2(n7374), 
        .Z(n1969) );
  OA22D0 U6030 ( .A1(n7375), .A2(prog_data[3]), .B1(\mem[168][3] ), .B2(n7374), 
        .Z(n1968) );
  OA22D0 U6031 ( .A1(n7375), .A2(prog_data[2]), .B1(\mem[168][2] ), .B2(n7374), 
        .Z(n1967) );
  OA22D0 U6032 ( .A1(n7375), .A2(prog_data[1]), .B1(\mem[168][1] ), .B2(n7374), 
        .Z(n1966) );
  OA22D0 U6033 ( .A1(n7375), .A2(prog_data[0]), .B1(\mem[168][0] ), .B2(n7374), 
        .Z(n1965) );
  NR2D0 U6034 ( .A1(n7555), .A2(n7388), .ZN(n7376) );
  INVD0 U6035 ( .I(n7376), .ZN(n7377) );
  OA22D0 U6036 ( .A1(n7377), .A2(prog_data[15]), .B1(\mem[169][15] ), .B2(
        n7376), .Z(n1964) );
  OA22D0 U6037 ( .A1(n7377), .A2(prog_data[14]), .B1(\mem[169][14] ), .B2(
        n7376), .Z(n1963) );
  OA22D0 U6038 ( .A1(n7377), .A2(prog_data[13]), .B1(\mem[169][13] ), .B2(
        n7376), .Z(n1962) );
  OA22D0 U6039 ( .A1(n7377), .A2(prog_data[12]), .B1(\mem[169][12] ), .B2(
        n7376), .Z(n1961) );
  OA22D0 U6040 ( .A1(n7377), .A2(prog_data[11]), .B1(\mem[169][11] ), .B2(
        n7376), .Z(n1960) );
  OA22D0 U6041 ( .A1(n7377), .A2(prog_data[10]), .B1(\mem[169][10] ), .B2(
        n7376), .Z(n1959) );
  OA22D0 U6042 ( .A1(n7377), .A2(prog_data[9]), .B1(\mem[169][9] ), .B2(n7376), 
        .Z(n1958) );
  OA22D0 U6043 ( .A1(n7377), .A2(prog_data[8]), .B1(\mem[169][8] ), .B2(n7376), 
        .Z(n1957) );
  OA22D0 U6044 ( .A1(n7377), .A2(prog_data[7]), .B1(\mem[169][7] ), .B2(n7376), 
        .Z(n1956) );
  OA22D0 U6045 ( .A1(n7377), .A2(prog_data[6]), .B1(\mem[169][6] ), .B2(n7376), 
        .Z(n1955) );
  OA22D0 U6046 ( .A1(n7377), .A2(prog_data[5]), .B1(\mem[169][5] ), .B2(n7376), 
        .Z(n1954) );
  OA22D0 U6047 ( .A1(n7377), .A2(prog_data[4]), .B1(\mem[169][4] ), .B2(n7376), 
        .Z(n1953) );
  OA22D0 U6048 ( .A1(n7377), .A2(prog_data[3]), .B1(\mem[169][3] ), .B2(n7376), 
        .Z(n1952) );
  OA22D0 U6049 ( .A1(n7377), .A2(prog_data[2]), .B1(\mem[169][2] ), .B2(n7376), 
        .Z(n1951) );
  OA22D0 U6050 ( .A1(n7377), .A2(prog_data[1]), .B1(\mem[169][1] ), .B2(n7376), 
        .Z(n1950) );
  OA22D0 U6051 ( .A1(n7377), .A2(prog_data[0]), .B1(\mem[169][0] ), .B2(n7376), 
        .Z(n1949) );
  NR2D0 U6052 ( .A1(n7558), .A2(n7388), .ZN(n7378) );
  INVD0 U6053 ( .I(n7378), .ZN(n7379) );
  OA22D0 U6054 ( .A1(n7379), .A2(prog_data[15]), .B1(\mem[170][15] ), .B2(
        n7378), .Z(n1948) );
  OA22D0 U6055 ( .A1(n7379), .A2(prog_data[14]), .B1(\mem[170][14] ), .B2(
        n7378), .Z(n1947) );
  OA22D0 U6056 ( .A1(n7379), .A2(prog_data[13]), .B1(\mem[170][13] ), .B2(
        n7378), .Z(n1946) );
  OA22D0 U6057 ( .A1(n7379), .A2(prog_data[12]), .B1(\mem[170][12] ), .B2(
        n7378), .Z(n1945) );
  OA22D0 U6058 ( .A1(n7379), .A2(prog_data[11]), .B1(\mem[170][11] ), .B2(
        n7378), .Z(n1944) );
  OA22D0 U6059 ( .A1(n7379), .A2(prog_data[10]), .B1(\mem[170][10] ), .B2(
        n7378), .Z(n1943) );
  OA22D0 U6060 ( .A1(n7379), .A2(prog_data[9]), .B1(\mem[170][9] ), .B2(n7378), 
        .Z(n1942) );
  OA22D0 U6061 ( .A1(n7379), .A2(prog_data[8]), .B1(\mem[170][8] ), .B2(n7378), 
        .Z(n1941) );
  OA22D0 U6062 ( .A1(n7379), .A2(prog_data[7]), .B1(\mem[170][7] ), .B2(n7378), 
        .Z(n1940) );
  OA22D0 U6063 ( .A1(n7379), .A2(prog_data[6]), .B1(\mem[170][6] ), .B2(n7378), 
        .Z(n1939) );
  OA22D0 U6064 ( .A1(n7379), .A2(prog_data[5]), .B1(\mem[170][5] ), .B2(n7378), 
        .Z(n1938) );
  OA22D0 U6065 ( .A1(n7379), .A2(prog_data[4]), .B1(\mem[170][4] ), .B2(n7378), 
        .Z(n1937) );
  OA22D0 U6066 ( .A1(n7379), .A2(prog_data[3]), .B1(\mem[170][3] ), .B2(n7378), 
        .Z(n1936) );
  OA22D0 U6067 ( .A1(n7379), .A2(prog_data[2]), .B1(\mem[170][2] ), .B2(n7378), 
        .Z(n1935) );
  OA22D0 U6068 ( .A1(n7379), .A2(prog_data[1]), .B1(\mem[170][1] ), .B2(n7378), 
        .Z(n1934) );
  OA22D0 U6069 ( .A1(n7379), .A2(prog_data[0]), .B1(\mem[170][0] ), .B2(n7378), 
        .Z(n1933) );
  NR2D0 U6070 ( .A1(n7561), .A2(n7388), .ZN(n7380) );
  INVD0 U6071 ( .I(n7380), .ZN(n7381) );
  OA22D0 U6072 ( .A1(n7381), .A2(prog_data[15]), .B1(\mem[171][15] ), .B2(
        n7380), .Z(n1932) );
  OA22D0 U6073 ( .A1(n7381), .A2(prog_data[14]), .B1(\mem[171][14] ), .B2(
        n7380), .Z(n1931) );
  OA22D0 U6074 ( .A1(n7381), .A2(prog_data[13]), .B1(\mem[171][13] ), .B2(
        n7380), .Z(n1930) );
  OA22D0 U6075 ( .A1(n7381), .A2(prog_data[12]), .B1(\mem[171][12] ), .B2(
        n7380), .Z(n1929) );
  OA22D0 U6076 ( .A1(n7381), .A2(prog_data[11]), .B1(\mem[171][11] ), .B2(
        n7380), .Z(n1928) );
  OA22D0 U6077 ( .A1(n7381), .A2(prog_data[10]), .B1(\mem[171][10] ), .B2(
        n7380), .Z(n1927) );
  OA22D0 U6078 ( .A1(n7381), .A2(prog_data[9]), .B1(\mem[171][9] ), .B2(n7380), 
        .Z(n1926) );
  OA22D0 U6079 ( .A1(n7381), .A2(prog_data[8]), .B1(\mem[171][8] ), .B2(n7380), 
        .Z(n1925) );
  OA22D0 U6080 ( .A1(n7381), .A2(prog_data[7]), .B1(\mem[171][7] ), .B2(n7380), 
        .Z(n1924) );
  OA22D0 U6081 ( .A1(n7381), .A2(prog_data[6]), .B1(\mem[171][6] ), .B2(n7380), 
        .Z(n1923) );
  OA22D0 U6082 ( .A1(n7381), .A2(prog_data[5]), .B1(\mem[171][5] ), .B2(n7380), 
        .Z(n1922) );
  OA22D0 U6083 ( .A1(n7381), .A2(prog_data[4]), .B1(\mem[171][4] ), .B2(n7380), 
        .Z(n1921) );
  OA22D0 U6084 ( .A1(n7381), .A2(prog_data[3]), .B1(\mem[171][3] ), .B2(n7380), 
        .Z(n1920) );
  OA22D0 U6085 ( .A1(n7381), .A2(prog_data[2]), .B1(\mem[171][2] ), .B2(n7380), 
        .Z(n1919) );
  OA22D0 U6086 ( .A1(n7381), .A2(prog_data[1]), .B1(\mem[171][1] ), .B2(n7380), 
        .Z(n1918) );
  OA22D0 U6087 ( .A1(n7381), .A2(prog_data[0]), .B1(\mem[171][0] ), .B2(n7380), 
        .Z(n1917) );
  NR2D0 U6088 ( .A1(n7564), .A2(n7388), .ZN(n7382) );
  INVD0 U6089 ( .I(n7382), .ZN(n7383) );
  OA22D0 U6090 ( .A1(n7383), .A2(prog_data[15]), .B1(\mem[172][15] ), .B2(
        n7382), .Z(n1916) );
  OA22D0 U6091 ( .A1(n7383), .A2(prog_data[14]), .B1(\mem[172][14] ), .B2(
        n7382), .Z(n1915) );
  OA22D0 U6092 ( .A1(n7383), .A2(prog_data[13]), .B1(\mem[172][13] ), .B2(
        n7382), .Z(n1914) );
  OA22D0 U6093 ( .A1(n7383), .A2(prog_data[12]), .B1(\mem[172][12] ), .B2(
        n7382), .Z(n1913) );
  OA22D0 U6094 ( .A1(n7383), .A2(prog_data[11]), .B1(\mem[172][11] ), .B2(
        n7382), .Z(n1912) );
  OA22D0 U6095 ( .A1(n7383), .A2(prog_data[10]), .B1(\mem[172][10] ), .B2(
        n7382), .Z(n1911) );
  OA22D0 U6096 ( .A1(n7383), .A2(prog_data[9]), .B1(\mem[172][9] ), .B2(n7382), 
        .Z(n1910) );
  OA22D0 U6097 ( .A1(n7383), .A2(prog_data[8]), .B1(\mem[172][8] ), .B2(n7382), 
        .Z(n1909) );
  OA22D0 U6098 ( .A1(n7383), .A2(prog_data[7]), .B1(\mem[172][7] ), .B2(n7382), 
        .Z(n1908) );
  OA22D0 U6099 ( .A1(n7383), .A2(prog_data[6]), .B1(\mem[172][6] ), .B2(n7382), 
        .Z(n1907) );
  OA22D0 U6100 ( .A1(n7383), .A2(prog_data[5]), .B1(\mem[172][5] ), .B2(n7382), 
        .Z(n1906) );
  OA22D0 U6101 ( .A1(n7383), .A2(prog_data[4]), .B1(\mem[172][4] ), .B2(n7382), 
        .Z(n1905) );
  OA22D0 U6102 ( .A1(n7383), .A2(prog_data[3]), .B1(\mem[172][3] ), .B2(n7382), 
        .Z(n1904) );
  OA22D0 U6103 ( .A1(n7383), .A2(prog_data[2]), .B1(\mem[172][2] ), .B2(n7382), 
        .Z(n1903) );
  OA22D0 U6104 ( .A1(n7383), .A2(prog_data[1]), .B1(\mem[172][1] ), .B2(n7382), 
        .Z(n1902) );
  OA22D0 U6105 ( .A1(n7383), .A2(prog_data[0]), .B1(\mem[172][0] ), .B2(n7382), 
        .Z(n1901) );
  NR2D0 U6106 ( .A1(n7567), .A2(n7388), .ZN(n7384) );
  INVD0 U6107 ( .I(n7384), .ZN(n7385) );
  OA22D0 U6108 ( .A1(n7385), .A2(prog_data[15]), .B1(\mem[173][15] ), .B2(
        n7384), .Z(n1900) );
  OA22D0 U6109 ( .A1(n7385), .A2(prog_data[14]), .B1(\mem[173][14] ), .B2(
        n7384), .Z(n1899) );
  OA22D0 U6110 ( .A1(n7385), .A2(prog_data[13]), .B1(\mem[173][13] ), .B2(
        n7384), .Z(n1898) );
  OA22D0 U6111 ( .A1(n7385), .A2(prog_data[12]), .B1(\mem[173][12] ), .B2(
        n7384), .Z(n1897) );
  OA22D0 U6112 ( .A1(n7385), .A2(prog_data[11]), .B1(\mem[173][11] ), .B2(
        n7384), .Z(n1896) );
  OA22D0 U6113 ( .A1(n7385), .A2(prog_data[10]), .B1(\mem[173][10] ), .B2(
        n7384), .Z(n1895) );
  OA22D0 U6114 ( .A1(n7385), .A2(prog_data[9]), .B1(\mem[173][9] ), .B2(n7384), 
        .Z(n1894) );
  OA22D0 U6115 ( .A1(n7385), .A2(prog_data[8]), .B1(\mem[173][8] ), .B2(n7384), 
        .Z(n1893) );
  OA22D0 U6116 ( .A1(n7385), .A2(prog_data[7]), .B1(\mem[173][7] ), .B2(n7384), 
        .Z(n1892) );
  OA22D0 U6117 ( .A1(n7385), .A2(prog_data[6]), .B1(\mem[173][6] ), .B2(n7384), 
        .Z(n1891) );
  OA22D0 U6118 ( .A1(n7385), .A2(prog_data[5]), .B1(\mem[173][5] ), .B2(n7384), 
        .Z(n1890) );
  OA22D0 U6119 ( .A1(n7385), .A2(prog_data[4]), .B1(\mem[173][4] ), .B2(n7384), 
        .Z(n1889) );
  OA22D0 U6120 ( .A1(n7385), .A2(prog_data[3]), .B1(\mem[173][3] ), .B2(n7384), 
        .Z(n1888) );
  OA22D0 U6121 ( .A1(n7385), .A2(prog_data[2]), .B1(\mem[173][2] ), .B2(n7384), 
        .Z(n1887) );
  OA22D0 U6122 ( .A1(n7385), .A2(prog_data[1]), .B1(\mem[173][1] ), .B2(n7384), 
        .Z(n1886) );
  OA22D0 U6123 ( .A1(n7385), .A2(prog_data[0]), .B1(\mem[173][0] ), .B2(n7384), 
        .Z(n1885) );
  NR2D0 U6124 ( .A1(n7570), .A2(n7388), .ZN(n7386) );
  OA22D0 U6125 ( .A1(n7387), .A2(prog_data[15]), .B1(\mem[174][15] ), .B2(
        n7386), .Z(n1884) );
  OA22D0 U6126 ( .A1(n7387), .A2(prog_data[14]), .B1(\mem[174][14] ), .B2(
        n7386), .Z(n1883) );
  OA22D0 U6127 ( .A1(n7387), .A2(prog_data[13]), .B1(\mem[174][13] ), .B2(
        n7386), .Z(n1882) );
  OA22D0 U6128 ( .A1(n7387), .A2(prog_data[12]), .B1(\mem[174][12] ), .B2(
        n7386), .Z(n1881) );
  OA22D0 U6129 ( .A1(n7387), .A2(prog_data[11]), .B1(\mem[174][11] ), .B2(
        n7386), .Z(n1880) );
  OA22D0 U6130 ( .A1(n7387), .A2(prog_data[10]), .B1(\mem[174][10] ), .B2(
        n7386), .Z(n1879) );
  OA22D0 U6131 ( .A1(n7387), .A2(prog_data[9]), .B1(\mem[174][9] ), .B2(n7386), 
        .Z(n1878) );
  OA22D0 U6132 ( .A1(n7387), .A2(prog_data[8]), .B1(\mem[174][8] ), .B2(n7386), 
        .Z(n1877) );
  OA22D0 U6133 ( .A1(n7387), .A2(prog_data[7]), .B1(\mem[174][7] ), .B2(n7386), 
        .Z(n1876) );
  OA22D0 U6134 ( .A1(n7387), .A2(prog_data[6]), .B1(\mem[174][6] ), .B2(n7386), 
        .Z(n1875) );
  OA22D0 U6135 ( .A1(n7387), .A2(prog_data[5]), .B1(\mem[174][5] ), .B2(n7386), 
        .Z(n1874) );
  OA22D0 U6136 ( .A1(n7387), .A2(prog_data[4]), .B1(\mem[174][4] ), .B2(n7386), 
        .Z(n1873) );
  OA22D0 U6137 ( .A1(n7387), .A2(prog_data[3]), .B1(\mem[174][3] ), .B2(n7386), 
        .Z(n1872) );
  OA22D0 U6138 ( .A1(n7387), .A2(prog_data[2]), .B1(\mem[174][2] ), .B2(n7386), 
        .Z(n1871) );
  OA22D0 U6139 ( .A1(n7387), .A2(prog_data[1]), .B1(\mem[174][1] ), .B2(n7386), 
        .Z(n1870) );
  OA22D0 U6140 ( .A1(n7387), .A2(prog_data[0]), .B1(\mem[174][0] ), .B2(n7386), 
        .Z(n1869) );
  NR2D0 U6141 ( .A1(n7574), .A2(n7388), .ZN(n7389) );
  INVD0 U6142 ( .I(n7389), .ZN(n7390) );
  OA22D0 U6143 ( .A1(n7390), .A2(prog_data[15]), .B1(\mem[175][15] ), .B2(
        n7389), .Z(n1868) );
  OA22D0 U6144 ( .A1(n7390), .A2(prog_data[14]), .B1(\mem[175][14] ), .B2(
        n7389), .Z(n1867) );
  OA22D0 U6145 ( .A1(n7390), .A2(prog_data[13]), .B1(\mem[175][13] ), .B2(
        n7389), .Z(n1866) );
  OA22D0 U6146 ( .A1(n7390), .A2(prog_data[12]), .B1(\mem[175][12] ), .B2(
        n7389), .Z(n1865) );
  OA22D0 U6147 ( .A1(n7390), .A2(prog_data[11]), .B1(\mem[175][11] ), .B2(
        n7389), .Z(n1864) );
  OA22D0 U6148 ( .A1(n7390), .A2(prog_data[10]), .B1(\mem[175][10] ), .B2(
        n7389), .Z(n1863) );
  OA22D0 U6149 ( .A1(n7390), .A2(prog_data[9]), .B1(\mem[175][9] ), .B2(n7389), 
        .Z(n1862) );
  OA22D0 U6150 ( .A1(n7390), .A2(prog_data[8]), .B1(\mem[175][8] ), .B2(n7389), 
        .Z(n1861) );
  OA22D0 U6151 ( .A1(n7390), .A2(prog_data[7]), .B1(\mem[175][7] ), .B2(n7389), 
        .Z(n1860) );
  OA22D0 U6152 ( .A1(n7390), .A2(prog_data[6]), .B1(\mem[175][6] ), .B2(n7389), 
        .Z(n1859) );
  OA22D0 U6153 ( .A1(n7390), .A2(prog_data[5]), .B1(\mem[175][5] ), .B2(n7389), 
        .Z(n1858) );
  OA22D0 U6154 ( .A1(n7390), .A2(prog_data[4]), .B1(\mem[175][4] ), .B2(n7389), 
        .Z(n1857) );
  OA22D0 U6155 ( .A1(n7390), .A2(prog_data[3]), .B1(\mem[175][3] ), .B2(n7389), 
        .Z(n1856) );
  OA22D0 U6156 ( .A1(n7390), .A2(prog_data[2]), .B1(\mem[175][2] ), .B2(n7389), 
        .Z(n1855) );
  OA22D0 U6157 ( .A1(n7390), .A2(prog_data[1]), .B1(\mem[175][1] ), .B2(n7389), 
        .Z(n1854) );
  OA22D0 U6158 ( .A1(n7390), .A2(prog_data[0]), .B1(\mem[175][0] ), .B2(n7389), 
        .Z(n1853) );
  CKND2D0 U6159 ( .A1(n7526), .A2(n7391), .ZN(n7422) );
  NR2D0 U6160 ( .A1(n7528), .A2(n7422), .ZN(n7392) );
  INVD0 U6161 ( .I(n7392), .ZN(n7393) );
  OA22D0 U6162 ( .A1(n7393), .A2(prog_data[15]), .B1(\mem[176][15] ), .B2(
        n7392), .Z(n1852) );
  OA22D0 U6163 ( .A1(n7393), .A2(prog_data[14]), .B1(\mem[176][14] ), .B2(
        n7392), .Z(n1851) );
  OA22D0 U6164 ( .A1(n7393), .A2(prog_data[13]), .B1(\mem[176][13] ), .B2(
        n7392), .Z(n1850) );
  OA22D0 U6165 ( .A1(n7393), .A2(prog_data[12]), .B1(\mem[176][12] ), .B2(
        n7392), .Z(n1849) );
  OA22D0 U6166 ( .A1(n7393), .A2(prog_data[11]), .B1(\mem[176][11] ), .B2(
        n7392), .Z(n1848) );
  OA22D0 U6167 ( .A1(n7393), .A2(prog_data[10]), .B1(\mem[176][10] ), .B2(
        n7392), .Z(n1847) );
  OA22D0 U6168 ( .A1(n7393), .A2(prog_data[9]), .B1(\mem[176][9] ), .B2(n7392), 
        .Z(n1846) );
  OA22D0 U6169 ( .A1(n7393), .A2(prog_data[8]), .B1(\mem[176][8] ), .B2(n7392), 
        .Z(n1845) );
  OA22D0 U6170 ( .A1(n7393), .A2(prog_data[7]), .B1(\mem[176][7] ), .B2(n7392), 
        .Z(n1844) );
  OA22D0 U6171 ( .A1(n7393), .A2(prog_data[6]), .B1(\mem[176][6] ), .B2(n7392), 
        .Z(n1843) );
  OA22D0 U6172 ( .A1(n7393), .A2(prog_data[5]), .B1(\mem[176][5] ), .B2(n7392), 
        .Z(n1842) );
  OA22D0 U6173 ( .A1(n7393), .A2(prog_data[4]), .B1(\mem[176][4] ), .B2(n7392), 
        .Z(n1841) );
  OA22D0 U6174 ( .A1(n7393), .A2(prog_data[3]), .B1(\mem[176][3] ), .B2(n7392), 
        .Z(n1840) );
  OA22D0 U6175 ( .A1(n7393), .A2(prog_data[2]), .B1(\mem[176][2] ), .B2(n7392), 
        .Z(n1839) );
  OA22D0 U6176 ( .A1(n7393), .A2(prog_data[1]), .B1(\mem[176][1] ), .B2(n7392), 
        .Z(n1838) );
  OA22D0 U6177 ( .A1(n7393), .A2(prog_data[0]), .B1(\mem[176][0] ), .B2(n7392), 
        .Z(n1837) );
  NR2D0 U6178 ( .A1(n7531), .A2(n7422), .ZN(n7394) );
  INVD0 U6179 ( .I(n7394), .ZN(n7395) );
  OA22D0 U6180 ( .A1(n7395), .A2(prog_data[15]), .B1(\mem[177][15] ), .B2(
        n7394), .Z(n1836) );
  OA22D0 U6181 ( .A1(n7395), .A2(prog_data[14]), .B1(\mem[177][14] ), .B2(
        n7394), .Z(n1835) );
  OA22D0 U6182 ( .A1(n7395), .A2(prog_data[13]), .B1(\mem[177][13] ), .B2(
        n7394), .Z(n1834) );
  OA22D0 U6183 ( .A1(n7395), .A2(prog_data[12]), .B1(\mem[177][12] ), .B2(
        n7394), .Z(n1833) );
  OA22D0 U6184 ( .A1(n7395), .A2(prog_data[11]), .B1(\mem[177][11] ), .B2(
        n7394), .Z(n1832) );
  OA22D0 U6185 ( .A1(n7395), .A2(prog_data[10]), .B1(\mem[177][10] ), .B2(
        n7394), .Z(n1831) );
  OA22D0 U6186 ( .A1(n7395), .A2(prog_data[9]), .B1(\mem[177][9] ), .B2(n7394), 
        .Z(n1830) );
  OA22D0 U6187 ( .A1(n7395), .A2(prog_data[8]), .B1(\mem[177][8] ), .B2(n7394), 
        .Z(n1829) );
  OA22D0 U6188 ( .A1(n7395), .A2(prog_data[7]), .B1(\mem[177][7] ), .B2(n7394), 
        .Z(n1828) );
  OA22D0 U6189 ( .A1(n7395), .A2(prog_data[6]), .B1(\mem[177][6] ), .B2(n7394), 
        .Z(n1827) );
  OA22D0 U6190 ( .A1(n7395), .A2(prog_data[5]), .B1(\mem[177][5] ), .B2(n7394), 
        .Z(n1826) );
  OA22D0 U6191 ( .A1(n7395), .A2(prog_data[4]), .B1(\mem[177][4] ), .B2(n7394), 
        .Z(n1825) );
  OA22D0 U6192 ( .A1(n7395), .A2(prog_data[3]), .B1(\mem[177][3] ), .B2(n7394), 
        .Z(n1824) );
  OA22D0 U6193 ( .A1(n7395), .A2(prog_data[2]), .B1(\mem[177][2] ), .B2(n7394), 
        .Z(n1823) );
  OA22D0 U6194 ( .A1(n7395), .A2(prog_data[1]), .B1(\mem[177][1] ), .B2(n7394), 
        .Z(n1822) );
  OA22D0 U6195 ( .A1(n7395), .A2(prog_data[0]), .B1(\mem[177][0] ), .B2(n7394), 
        .Z(n1821) );
  NR2D0 U6196 ( .A1(n7534), .A2(n7422), .ZN(n7396) );
  INVD0 U6197 ( .I(n7396), .ZN(n7397) );
  OA22D0 U6198 ( .A1(n7397), .A2(prog_data[15]), .B1(\mem[178][15] ), .B2(
        n7396), .Z(n1820) );
  OA22D0 U6199 ( .A1(n7397), .A2(prog_data[14]), .B1(\mem[178][14] ), .B2(
        n7396), .Z(n1819) );
  OA22D0 U6200 ( .A1(n7397), .A2(prog_data[13]), .B1(\mem[178][13] ), .B2(
        n7396), .Z(n1818) );
  OA22D0 U6201 ( .A1(n7397), .A2(prog_data[12]), .B1(\mem[178][12] ), .B2(
        n7396), .Z(n1817) );
  OA22D0 U6202 ( .A1(n7397), .A2(prog_data[11]), .B1(\mem[178][11] ), .B2(
        n7396), .Z(n1816) );
  OA22D0 U6203 ( .A1(n7397), .A2(prog_data[10]), .B1(\mem[178][10] ), .B2(
        n7396), .Z(n1815) );
  OA22D0 U6204 ( .A1(n7397), .A2(prog_data[9]), .B1(\mem[178][9] ), .B2(n7396), 
        .Z(n1814) );
  OA22D0 U6205 ( .A1(n7397), .A2(prog_data[8]), .B1(\mem[178][8] ), .B2(n7396), 
        .Z(n1813) );
  OA22D0 U6206 ( .A1(n7397), .A2(prog_data[7]), .B1(\mem[178][7] ), .B2(n7396), 
        .Z(n1812) );
  OA22D0 U6207 ( .A1(n7397), .A2(prog_data[6]), .B1(\mem[178][6] ), .B2(n7396), 
        .Z(n1811) );
  OA22D0 U6208 ( .A1(n7397), .A2(prog_data[5]), .B1(\mem[178][5] ), .B2(n7396), 
        .Z(n1810) );
  OA22D0 U6209 ( .A1(n7397), .A2(prog_data[4]), .B1(\mem[178][4] ), .B2(n7396), 
        .Z(n1809) );
  OA22D0 U6210 ( .A1(n7397), .A2(prog_data[3]), .B1(\mem[178][3] ), .B2(n7396), 
        .Z(n1808) );
  OA22D0 U6211 ( .A1(n7397), .A2(prog_data[2]), .B1(\mem[178][2] ), .B2(n7396), 
        .Z(n1807) );
  OA22D0 U6212 ( .A1(n7397), .A2(prog_data[1]), .B1(\mem[178][1] ), .B2(n7396), 
        .Z(n1806) );
  OA22D0 U6213 ( .A1(n7397), .A2(prog_data[0]), .B1(\mem[178][0] ), .B2(n7396), 
        .Z(n1805) );
  NR2D0 U6214 ( .A1(n7537), .A2(n7422), .ZN(n7398) );
  INVD0 U6215 ( .I(n7398), .ZN(n7399) );
  OA22D0 U6216 ( .A1(n7399), .A2(prog_data[15]), .B1(\mem[179][15] ), .B2(
        n7398), .Z(n1804) );
  OA22D0 U6217 ( .A1(n7399), .A2(prog_data[14]), .B1(\mem[179][14] ), .B2(
        n7398), .Z(n1803) );
  OA22D0 U6218 ( .A1(n7399), .A2(prog_data[13]), .B1(\mem[179][13] ), .B2(
        n7398), .Z(n1802) );
  OA22D0 U6219 ( .A1(n7399), .A2(prog_data[12]), .B1(\mem[179][12] ), .B2(
        n7398), .Z(n1801) );
  OA22D0 U6220 ( .A1(n7399), .A2(prog_data[11]), .B1(\mem[179][11] ), .B2(
        n7398), .Z(n1800) );
  OA22D0 U6221 ( .A1(n7399), .A2(prog_data[10]), .B1(\mem[179][10] ), .B2(
        n7398), .Z(n1799) );
  OA22D0 U6222 ( .A1(n7399), .A2(prog_data[9]), .B1(\mem[179][9] ), .B2(n7398), 
        .Z(n1798) );
  OA22D0 U6223 ( .A1(n7399), .A2(prog_data[8]), .B1(\mem[179][8] ), .B2(n7398), 
        .Z(n1797) );
  OA22D0 U6224 ( .A1(n7399), .A2(prog_data[7]), .B1(\mem[179][7] ), .B2(n7398), 
        .Z(n1796) );
  OA22D0 U6225 ( .A1(n7399), .A2(prog_data[6]), .B1(\mem[179][6] ), .B2(n7398), 
        .Z(n1795) );
  OA22D0 U6226 ( .A1(n7399), .A2(prog_data[5]), .B1(\mem[179][5] ), .B2(n7398), 
        .Z(n1794) );
  OA22D0 U6227 ( .A1(n7399), .A2(prog_data[4]), .B1(\mem[179][4] ), .B2(n7398), 
        .Z(n1793) );
  OA22D0 U6228 ( .A1(n7399), .A2(prog_data[3]), .B1(\mem[179][3] ), .B2(n7398), 
        .Z(n1792) );
  OA22D0 U6229 ( .A1(n7399), .A2(prog_data[2]), .B1(\mem[179][2] ), .B2(n7398), 
        .Z(n1791) );
  OA22D0 U6230 ( .A1(n7399), .A2(prog_data[1]), .B1(\mem[179][1] ), .B2(n7398), 
        .Z(n1790) );
  OA22D0 U6231 ( .A1(n7399), .A2(prog_data[0]), .B1(\mem[179][0] ), .B2(n7398), 
        .Z(n1789) );
  NR2D0 U6232 ( .A1(n7540), .A2(n7422), .ZN(n7400) );
  INVD0 U6233 ( .I(n7400), .ZN(n7401) );
  OA22D0 U6234 ( .A1(n7401), .A2(prog_data[15]), .B1(\mem[180][15] ), .B2(
        n7400), .Z(n1788) );
  OA22D0 U6235 ( .A1(n7401), .A2(prog_data[14]), .B1(\mem[180][14] ), .B2(
        n7400), .Z(n1787) );
  OA22D0 U6236 ( .A1(n7401), .A2(prog_data[13]), .B1(\mem[180][13] ), .B2(
        n7400), .Z(n1786) );
  OA22D0 U6237 ( .A1(n7401), .A2(prog_data[12]), .B1(\mem[180][12] ), .B2(
        n7400), .Z(n1785) );
  OA22D0 U6238 ( .A1(n7401), .A2(prog_data[11]), .B1(\mem[180][11] ), .B2(
        n7400), .Z(n1784) );
  OA22D0 U6239 ( .A1(n7401), .A2(prog_data[10]), .B1(\mem[180][10] ), .B2(
        n7400), .Z(n1783) );
  OA22D0 U6240 ( .A1(n7401), .A2(prog_data[9]), .B1(\mem[180][9] ), .B2(n7400), 
        .Z(n1782) );
  OA22D0 U6241 ( .A1(n7401), .A2(prog_data[8]), .B1(\mem[180][8] ), .B2(n7400), 
        .Z(n1781) );
  OA22D0 U6242 ( .A1(n7401), .A2(prog_data[7]), .B1(\mem[180][7] ), .B2(n7400), 
        .Z(n1780) );
  OA22D0 U6243 ( .A1(n7401), .A2(prog_data[6]), .B1(\mem[180][6] ), .B2(n7400), 
        .Z(n1779) );
  OA22D0 U6244 ( .A1(n7401), .A2(prog_data[5]), .B1(\mem[180][5] ), .B2(n7400), 
        .Z(n1778) );
  OA22D0 U6245 ( .A1(n7401), .A2(prog_data[4]), .B1(\mem[180][4] ), .B2(n7400), 
        .Z(n1777) );
  OA22D0 U6246 ( .A1(n7401), .A2(prog_data[3]), .B1(\mem[180][3] ), .B2(n7400), 
        .Z(n1776) );
  OA22D0 U6247 ( .A1(n7401), .A2(prog_data[2]), .B1(\mem[180][2] ), .B2(n7400), 
        .Z(n1775) );
  OA22D0 U6248 ( .A1(n7401), .A2(prog_data[1]), .B1(\mem[180][1] ), .B2(n7400), 
        .Z(n1774) );
  OA22D0 U6249 ( .A1(n7401), .A2(prog_data[0]), .B1(\mem[180][0] ), .B2(n7400), 
        .Z(n1773) );
  INVD0 U6250 ( .I(n7402), .ZN(n7403) );
  OA22D0 U6251 ( .A1(n7403), .A2(prog_data[15]), .B1(\mem[181][15] ), .B2(
        n7402), .Z(n1772) );
  OA22D0 U6252 ( .A1(n7403), .A2(prog_data[14]), .B1(\mem[181][14] ), .B2(
        n7402), .Z(n1771) );
  OA22D0 U6253 ( .A1(n7403), .A2(prog_data[13]), .B1(\mem[181][13] ), .B2(
        n7402), .Z(n1770) );
  OA22D0 U6254 ( .A1(n7403), .A2(prog_data[12]), .B1(\mem[181][12] ), .B2(
        n7402), .Z(n1769) );
  OA22D0 U6255 ( .A1(n7403), .A2(prog_data[11]), .B1(\mem[181][11] ), .B2(
        n7402), .Z(n1768) );
  OA22D0 U6256 ( .A1(n7403), .A2(prog_data[10]), .B1(\mem[181][10] ), .B2(
        n7402), .Z(n1767) );
  OA22D0 U6257 ( .A1(n7403), .A2(prog_data[9]), .B1(\mem[181][9] ), .B2(n7402), 
        .Z(n1766) );
  OA22D0 U6258 ( .A1(n7403), .A2(prog_data[8]), .B1(\mem[181][8] ), .B2(n7402), 
        .Z(n1765) );
  OA22D0 U6259 ( .A1(n7403), .A2(prog_data[7]), .B1(\mem[181][7] ), .B2(n7402), 
        .Z(n1764) );
  OA22D0 U6260 ( .A1(n7403), .A2(prog_data[6]), .B1(\mem[181][6] ), .B2(n7402), 
        .Z(n1763) );
  OA22D0 U6261 ( .A1(n7403), .A2(prog_data[5]), .B1(\mem[181][5] ), .B2(n7402), 
        .Z(n1762) );
  OA22D0 U6262 ( .A1(n7403), .A2(prog_data[4]), .B1(\mem[181][4] ), .B2(n7402), 
        .Z(n1761) );
  OA22D0 U6263 ( .A1(n7403), .A2(prog_data[3]), .B1(\mem[181][3] ), .B2(n7402), 
        .Z(n1760) );
  OA22D0 U6264 ( .A1(n7403), .A2(prog_data[2]), .B1(\mem[181][2] ), .B2(n7402), 
        .Z(n1759) );
  OA22D0 U6265 ( .A1(n7403), .A2(prog_data[1]), .B1(\mem[181][1] ), .B2(n7402), 
        .Z(n1758) );
  OA22D0 U6266 ( .A1(n7403), .A2(prog_data[0]), .B1(\mem[181][0] ), .B2(n7402), 
        .Z(n1757) );
  NR2D0 U6267 ( .A1(n7546), .A2(n7422), .ZN(n7404) );
  INVD0 U6268 ( .I(n7404), .ZN(n7405) );
  OA22D0 U6269 ( .A1(n7405), .A2(prog_data[15]), .B1(\mem[182][15] ), .B2(
        n7404), .Z(n1756) );
  OA22D0 U6270 ( .A1(n7405), .A2(prog_data[14]), .B1(\mem[182][14] ), .B2(
        n7404), .Z(n1755) );
  OA22D0 U6271 ( .A1(n7405), .A2(prog_data[13]), .B1(\mem[182][13] ), .B2(
        n7404), .Z(n1754) );
  OA22D0 U6272 ( .A1(n7405), .A2(prog_data[12]), .B1(\mem[182][12] ), .B2(
        n7404), .Z(n1753) );
  OA22D0 U6273 ( .A1(n7405), .A2(prog_data[11]), .B1(\mem[182][11] ), .B2(
        n7404), .Z(n1752) );
  OA22D0 U6274 ( .A1(n7405), .A2(prog_data[10]), .B1(\mem[182][10] ), .B2(
        n7404), .Z(n1751) );
  OA22D0 U6275 ( .A1(n7405), .A2(prog_data[9]), .B1(\mem[182][9] ), .B2(n7404), 
        .Z(n1750) );
  OA22D0 U6276 ( .A1(n7405), .A2(prog_data[8]), .B1(\mem[182][8] ), .B2(n7404), 
        .Z(n1749) );
  OA22D0 U6277 ( .A1(n7405), .A2(prog_data[7]), .B1(\mem[182][7] ), .B2(n7404), 
        .Z(n1748) );
  OA22D0 U6278 ( .A1(n7405), .A2(prog_data[6]), .B1(\mem[182][6] ), .B2(n7404), 
        .Z(n1747) );
  OA22D0 U6279 ( .A1(n7405), .A2(prog_data[5]), .B1(\mem[182][5] ), .B2(n7404), 
        .Z(n1746) );
  OA22D0 U6280 ( .A1(n7405), .A2(prog_data[4]), .B1(\mem[182][4] ), .B2(n7404), 
        .Z(n1745) );
  OA22D0 U6281 ( .A1(n7405), .A2(prog_data[3]), .B1(\mem[182][3] ), .B2(n7404), 
        .Z(n1744) );
  OA22D0 U6282 ( .A1(n7405), .A2(prog_data[2]), .B1(\mem[182][2] ), .B2(n7404), 
        .Z(n1743) );
  OA22D0 U6283 ( .A1(n7405), .A2(prog_data[1]), .B1(\mem[182][1] ), .B2(n7404), 
        .Z(n1742) );
  OA22D0 U6284 ( .A1(n7405), .A2(prog_data[0]), .B1(\mem[182][0] ), .B2(n7404), 
        .Z(n1741) );
  NR2D0 U6285 ( .A1(n7549), .A2(n7422), .ZN(n7406) );
  INVD0 U6286 ( .I(n7406), .ZN(n7407) );
  OA22D0 U6287 ( .A1(n7407), .A2(prog_data[15]), .B1(\mem[183][15] ), .B2(
        n7406), .Z(n1740) );
  OA22D0 U6288 ( .A1(n7407), .A2(prog_data[14]), .B1(\mem[183][14] ), .B2(
        n7406), .Z(n1739) );
  OA22D0 U6289 ( .A1(n7407), .A2(prog_data[13]), .B1(\mem[183][13] ), .B2(
        n7406), .Z(n1738) );
  OA22D0 U6290 ( .A1(n7407), .A2(prog_data[12]), .B1(\mem[183][12] ), .B2(
        n7406), .Z(n1737) );
  OA22D0 U6291 ( .A1(n7407), .A2(prog_data[11]), .B1(\mem[183][11] ), .B2(
        n7406), .Z(n1736) );
  OA22D0 U6292 ( .A1(n7407), .A2(prog_data[10]), .B1(\mem[183][10] ), .B2(
        n7406), .Z(n1735) );
  OA22D0 U6293 ( .A1(n7407), .A2(prog_data[9]), .B1(\mem[183][9] ), .B2(n7406), 
        .Z(n1734) );
  OA22D0 U6294 ( .A1(n7407), .A2(prog_data[8]), .B1(\mem[183][8] ), .B2(n7406), 
        .Z(n1733) );
  OA22D0 U6295 ( .A1(n7407), .A2(prog_data[7]), .B1(\mem[183][7] ), .B2(n7406), 
        .Z(n1732) );
  OA22D0 U6296 ( .A1(n7407), .A2(prog_data[6]), .B1(\mem[183][6] ), .B2(n7406), 
        .Z(n1731) );
  OA22D0 U6297 ( .A1(n7407), .A2(prog_data[5]), .B1(\mem[183][5] ), .B2(n7406), 
        .Z(n1730) );
  OA22D0 U6298 ( .A1(n7407), .A2(prog_data[4]), .B1(\mem[183][4] ), .B2(n7406), 
        .Z(n1729) );
  OA22D0 U6299 ( .A1(n7407), .A2(prog_data[3]), .B1(\mem[183][3] ), .B2(n7406), 
        .Z(n1728) );
  OA22D0 U6300 ( .A1(n7407), .A2(prog_data[2]), .B1(\mem[183][2] ), .B2(n7406), 
        .Z(n1727) );
  OA22D0 U6301 ( .A1(n7407), .A2(prog_data[1]), .B1(\mem[183][1] ), .B2(n7406), 
        .Z(n1726) );
  OA22D0 U6302 ( .A1(n7407), .A2(prog_data[0]), .B1(\mem[183][0] ), .B2(n7406), 
        .Z(n1725) );
  NR2D0 U6303 ( .A1(n7552), .A2(n7422), .ZN(n7408) );
  INVD0 U6304 ( .I(n7408), .ZN(n7409) );
  OA22D0 U6305 ( .A1(n7409), .A2(prog_data[15]), .B1(\mem[184][15] ), .B2(
        n7408), .Z(n1724) );
  OA22D0 U6306 ( .A1(n7409), .A2(prog_data[14]), .B1(\mem[184][14] ), .B2(
        n7408), .Z(n1723) );
  OA22D0 U6307 ( .A1(n7409), .A2(prog_data[13]), .B1(\mem[184][13] ), .B2(
        n7408), .Z(n1722) );
  OA22D0 U6308 ( .A1(n7409), .A2(prog_data[12]), .B1(\mem[184][12] ), .B2(
        n7408), .Z(n1721) );
  OA22D0 U6309 ( .A1(n7409), .A2(prog_data[11]), .B1(\mem[184][11] ), .B2(
        n7408), .Z(n1720) );
  OA22D0 U6310 ( .A1(n7409), .A2(prog_data[10]), .B1(\mem[184][10] ), .B2(
        n7408), .Z(n1719) );
  OA22D0 U6311 ( .A1(n7409), .A2(prog_data[9]), .B1(\mem[184][9] ), .B2(n7408), 
        .Z(n1718) );
  OA22D0 U6312 ( .A1(n7409), .A2(prog_data[8]), .B1(\mem[184][8] ), .B2(n7408), 
        .Z(n1717) );
  OA22D0 U6313 ( .A1(n7409), .A2(prog_data[7]), .B1(\mem[184][7] ), .B2(n7408), 
        .Z(n1716) );
  OA22D0 U6314 ( .A1(n7409), .A2(prog_data[6]), .B1(\mem[184][6] ), .B2(n7408), 
        .Z(n1715) );
  OA22D0 U6315 ( .A1(n7409), .A2(prog_data[5]), .B1(\mem[184][5] ), .B2(n7408), 
        .Z(n1714) );
  OA22D0 U6316 ( .A1(n7409), .A2(prog_data[4]), .B1(\mem[184][4] ), .B2(n7408), 
        .Z(n1713) );
  OA22D0 U6317 ( .A1(n7409), .A2(prog_data[3]), .B1(\mem[184][3] ), .B2(n7408), 
        .Z(n1712) );
  OA22D0 U6318 ( .A1(n7409), .A2(prog_data[2]), .B1(\mem[184][2] ), .B2(n7408), 
        .Z(n1711) );
  OA22D0 U6319 ( .A1(n7409), .A2(prog_data[1]), .B1(\mem[184][1] ), .B2(n7408), 
        .Z(n1710) );
  OA22D0 U6320 ( .A1(n7409), .A2(prog_data[0]), .B1(\mem[184][0] ), .B2(n7408), 
        .Z(n1709) );
  NR2D0 U6321 ( .A1(n7555), .A2(n7422), .ZN(n7410) );
  INVD0 U6322 ( .I(n7410), .ZN(n7411) );
  OA22D0 U6323 ( .A1(n7411), .A2(prog_data[15]), .B1(\mem[185][15] ), .B2(
        n7410), .Z(n1708) );
  OA22D0 U6324 ( .A1(n7411), .A2(prog_data[14]), .B1(\mem[185][14] ), .B2(
        n7410), .Z(n1707) );
  OA22D0 U6325 ( .A1(n7411), .A2(prog_data[13]), .B1(\mem[185][13] ), .B2(
        n7410), .Z(n1706) );
  OA22D0 U6326 ( .A1(n7411), .A2(prog_data[12]), .B1(\mem[185][12] ), .B2(
        n7410), .Z(n1705) );
  OA22D0 U6327 ( .A1(n7411), .A2(prog_data[11]), .B1(\mem[185][11] ), .B2(
        n7410), .Z(n1704) );
  OA22D0 U6328 ( .A1(n7411), .A2(prog_data[10]), .B1(\mem[185][10] ), .B2(
        n7410), .Z(n1703) );
  OA22D0 U6329 ( .A1(n7411), .A2(prog_data[9]), .B1(\mem[185][9] ), .B2(n7410), 
        .Z(n1702) );
  OA22D0 U6330 ( .A1(n7411), .A2(prog_data[8]), .B1(\mem[185][8] ), .B2(n7410), 
        .Z(n1701) );
  OA22D0 U6331 ( .A1(n7411), .A2(prog_data[7]), .B1(\mem[185][7] ), .B2(n7410), 
        .Z(n1700) );
  OA22D0 U6332 ( .A1(n7411), .A2(prog_data[6]), .B1(\mem[185][6] ), .B2(n7410), 
        .Z(n1699) );
  OA22D0 U6333 ( .A1(n7411), .A2(prog_data[5]), .B1(\mem[185][5] ), .B2(n7410), 
        .Z(n1698) );
  OA22D0 U6334 ( .A1(n7411), .A2(prog_data[4]), .B1(\mem[185][4] ), .B2(n7410), 
        .Z(n1697) );
  OA22D0 U6335 ( .A1(n7411), .A2(prog_data[3]), .B1(\mem[185][3] ), .B2(n7410), 
        .Z(n1696) );
  OA22D0 U6336 ( .A1(n7411), .A2(prog_data[2]), .B1(\mem[185][2] ), .B2(n7410), 
        .Z(n1695) );
  OA22D0 U6337 ( .A1(n7411), .A2(prog_data[1]), .B1(\mem[185][1] ), .B2(n7410), 
        .Z(n1694) );
  OA22D0 U6338 ( .A1(n7411), .A2(prog_data[0]), .B1(\mem[185][0] ), .B2(n7410), 
        .Z(n1693) );
  NR2D0 U6339 ( .A1(n7558), .A2(n7422), .ZN(n7412) );
  INVD0 U6340 ( .I(n7412), .ZN(n7413) );
  OA22D0 U6341 ( .A1(n7413), .A2(prog_data[15]), .B1(\mem[186][15] ), .B2(
        n7412), .Z(n1692) );
  OA22D0 U6342 ( .A1(n7413), .A2(prog_data[14]), .B1(\mem[186][14] ), .B2(
        n7412), .Z(n1691) );
  OA22D0 U6343 ( .A1(n7413), .A2(prog_data[13]), .B1(\mem[186][13] ), .B2(
        n7412), .Z(n1690) );
  OA22D0 U6344 ( .A1(n7413), .A2(prog_data[12]), .B1(\mem[186][12] ), .B2(
        n7412), .Z(n1689) );
  OA22D0 U6345 ( .A1(n7413), .A2(prog_data[11]), .B1(\mem[186][11] ), .B2(
        n7412), .Z(n1688) );
  OA22D0 U6346 ( .A1(n7413), .A2(prog_data[10]), .B1(\mem[186][10] ), .B2(
        n7412), .Z(n1687) );
  OA22D0 U6347 ( .A1(n7413), .A2(prog_data[9]), .B1(\mem[186][9] ), .B2(n7412), 
        .Z(n1686) );
  OA22D0 U6348 ( .A1(n7413), .A2(prog_data[8]), .B1(\mem[186][8] ), .B2(n7412), 
        .Z(n1685) );
  OA22D0 U6349 ( .A1(n7413), .A2(prog_data[7]), .B1(\mem[186][7] ), .B2(n7412), 
        .Z(n1684) );
  OA22D0 U6350 ( .A1(n7413), .A2(prog_data[6]), .B1(\mem[186][6] ), .B2(n7412), 
        .Z(n1683) );
  OA22D0 U6351 ( .A1(n7413), .A2(prog_data[5]), .B1(\mem[186][5] ), .B2(n7412), 
        .Z(n1682) );
  OA22D0 U6352 ( .A1(n7413), .A2(prog_data[4]), .B1(\mem[186][4] ), .B2(n7412), 
        .Z(n1681) );
  OA22D0 U6353 ( .A1(n7413), .A2(prog_data[3]), .B1(\mem[186][3] ), .B2(n7412), 
        .Z(n1680) );
  OA22D0 U6354 ( .A1(n7413), .A2(prog_data[2]), .B1(\mem[186][2] ), .B2(n7412), 
        .Z(n1679) );
  OA22D0 U6355 ( .A1(n7413), .A2(prog_data[1]), .B1(\mem[186][1] ), .B2(n7412), 
        .Z(n1678) );
  OA22D0 U6356 ( .A1(n7413), .A2(prog_data[0]), .B1(\mem[186][0] ), .B2(n7412), 
        .Z(n1677) );
  NR2D0 U6357 ( .A1(n7561), .A2(n7422), .ZN(n7414) );
  INVD0 U6358 ( .I(n7414), .ZN(n7415) );
  OA22D0 U6359 ( .A1(n7415), .A2(prog_data[15]), .B1(\mem[187][15] ), .B2(
        n7414), .Z(n1676) );
  OA22D0 U6360 ( .A1(n7415), .A2(prog_data[14]), .B1(\mem[187][14] ), .B2(
        n7414), .Z(n1675) );
  OA22D0 U6361 ( .A1(n7415), .A2(prog_data[13]), .B1(\mem[187][13] ), .B2(
        n7414), .Z(n1674) );
  OA22D0 U6362 ( .A1(n7415), .A2(prog_data[12]), .B1(\mem[187][12] ), .B2(
        n7414), .Z(n1673) );
  OA22D0 U6363 ( .A1(n7415), .A2(prog_data[11]), .B1(\mem[187][11] ), .B2(
        n7414), .Z(n1672) );
  OA22D0 U6364 ( .A1(n7415), .A2(prog_data[10]), .B1(\mem[187][10] ), .B2(
        n7414), .Z(n1671) );
  OA22D0 U6365 ( .A1(n7415), .A2(prog_data[9]), .B1(\mem[187][9] ), .B2(n7414), 
        .Z(n1670) );
  OA22D0 U6366 ( .A1(n7415), .A2(prog_data[8]), .B1(\mem[187][8] ), .B2(n7414), 
        .Z(n1669) );
  OA22D0 U6367 ( .A1(n7415), .A2(prog_data[7]), .B1(\mem[187][7] ), .B2(n7414), 
        .Z(n1668) );
  OA22D0 U6368 ( .A1(n7415), .A2(prog_data[6]), .B1(\mem[187][6] ), .B2(n7414), 
        .Z(n1667) );
  OA22D0 U6369 ( .A1(n7415), .A2(prog_data[5]), .B1(\mem[187][5] ), .B2(n7414), 
        .Z(n1666) );
  OA22D0 U6370 ( .A1(n7415), .A2(prog_data[4]), .B1(\mem[187][4] ), .B2(n7414), 
        .Z(n1665) );
  OA22D0 U6371 ( .A1(n7415), .A2(prog_data[3]), .B1(\mem[187][3] ), .B2(n7414), 
        .Z(n1664) );
  OA22D0 U6372 ( .A1(n7415), .A2(prog_data[2]), .B1(\mem[187][2] ), .B2(n7414), 
        .Z(n1663) );
  OA22D0 U6373 ( .A1(n7415), .A2(prog_data[1]), .B1(\mem[187][1] ), .B2(n7414), 
        .Z(n1662) );
  OA22D0 U6374 ( .A1(n7415), .A2(prog_data[0]), .B1(\mem[187][0] ), .B2(n7414), 
        .Z(n1661) );
  NR2D0 U6375 ( .A1(n7564), .A2(n7422), .ZN(n7416) );
  INVD0 U6376 ( .I(n7416), .ZN(n7417) );
  OA22D0 U6377 ( .A1(n7417), .A2(prog_data[15]), .B1(\mem[188][15] ), .B2(
        n7416), .Z(n1660) );
  OA22D0 U6378 ( .A1(n7417), .A2(prog_data[14]), .B1(\mem[188][14] ), .B2(
        n7416), .Z(n1659) );
  OA22D0 U6379 ( .A1(n7417), .A2(prog_data[13]), .B1(\mem[188][13] ), .B2(
        n7416), .Z(n1658) );
  OA22D0 U6380 ( .A1(n7417), .A2(prog_data[12]), .B1(\mem[188][12] ), .B2(
        n7416), .Z(n1657) );
  OA22D0 U6381 ( .A1(n7417), .A2(prog_data[11]), .B1(\mem[188][11] ), .B2(
        n7416), .Z(n1656) );
  OA22D0 U6382 ( .A1(n7417), .A2(prog_data[10]), .B1(\mem[188][10] ), .B2(
        n7416), .Z(n1655) );
  OA22D0 U6383 ( .A1(n7417), .A2(prog_data[9]), .B1(\mem[188][9] ), .B2(n7416), 
        .Z(n1654) );
  OA22D0 U6384 ( .A1(n7417), .A2(prog_data[8]), .B1(\mem[188][8] ), .B2(n7416), 
        .Z(n1653) );
  OA22D0 U6385 ( .A1(n7417), .A2(prog_data[7]), .B1(\mem[188][7] ), .B2(n7416), 
        .Z(n1652) );
  OA22D0 U6386 ( .A1(n7417), .A2(prog_data[6]), .B1(\mem[188][6] ), .B2(n7416), 
        .Z(n1651) );
  OA22D0 U6387 ( .A1(n7417), .A2(prog_data[5]), .B1(\mem[188][5] ), .B2(n7416), 
        .Z(n1650) );
  OA22D0 U6388 ( .A1(n7417), .A2(prog_data[4]), .B1(\mem[188][4] ), .B2(n7416), 
        .Z(n1649) );
  OA22D0 U6389 ( .A1(n7417), .A2(prog_data[3]), .B1(\mem[188][3] ), .B2(n7416), 
        .Z(n1648) );
  OA22D0 U6390 ( .A1(n7417), .A2(prog_data[2]), .B1(\mem[188][2] ), .B2(n7416), 
        .Z(n1647) );
  OA22D0 U6391 ( .A1(n7417), .A2(prog_data[1]), .B1(\mem[188][1] ), .B2(n7416), 
        .Z(n1646) );
  OA22D0 U6392 ( .A1(n7417), .A2(prog_data[0]), .B1(\mem[188][0] ), .B2(n7416), 
        .Z(n1645) );
  NR2D0 U6393 ( .A1(n7567), .A2(n7422), .ZN(n7418) );
  OA22D0 U6394 ( .A1(n7419), .A2(prog_data[15]), .B1(\mem[189][15] ), .B2(
        n7418), .Z(n1644) );
  OA22D0 U6395 ( .A1(n7419), .A2(prog_data[14]), .B1(\mem[189][14] ), .B2(
        n7418), .Z(n1643) );
  OA22D0 U6396 ( .A1(n7419), .A2(prog_data[13]), .B1(\mem[189][13] ), .B2(
        n7418), .Z(n1642) );
  OA22D0 U6397 ( .A1(n7419), .A2(prog_data[12]), .B1(\mem[189][12] ), .B2(
        n7418), .Z(n1641) );
  OA22D0 U6398 ( .A1(n7419), .A2(prog_data[11]), .B1(\mem[189][11] ), .B2(
        n7418), .Z(n1640) );
  OA22D0 U6399 ( .A1(n7419), .A2(prog_data[10]), .B1(\mem[189][10] ), .B2(
        n7418), .Z(n1639) );
  OA22D0 U6400 ( .A1(n7419), .A2(prog_data[9]), .B1(\mem[189][9] ), .B2(n7418), 
        .Z(n1638) );
  OA22D0 U6401 ( .A1(n7419), .A2(prog_data[8]), .B1(\mem[189][8] ), .B2(n7418), 
        .Z(n1637) );
  OA22D0 U6402 ( .A1(n7419), .A2(prog_data[7]), .B1(\mem[189][7] ), .B2(n7418), 
        .Z(n1636) );
  OA22D0 U6403 ( .A1(n7419), .A2(prog_data[6]), .B1(\mem[189][6] ), .B2(n7418), 
        .Z(n1635) );
  OA22D0 U6404 ( .A1(n7419), .A2(prog_data[5]), .B1(\mem[189][5] ), .B2(n7418), 
        .Z(n1634) );
  OA22D0 U6405 ( .A1(n7419), .A2(prog_data[4]), .B1(\mem[189][4] ), .B2(n7418), 
        .Z(n1633) );
  OA22D0 U6406 ( .A1(n7419), .A2(prog_data[3]), .B1(\mem[189][3] ), .B2(n7418), 
        .Z(n1632) );
  OA22D0 U6407 ( .A1(n7419), .A2(prog_data[2]), .B1(\mem[189][2] ), .B2(n7418), 
        .Z(n1631) );
  OA22D0 U6408 ( .A1(n7419), .A2(prog_data[1]), .B1(\mem[189][1] ), .B2(n7418), 
        .Z(n1630) );
  OA22D0 U6409 ( .A1(n7419), .A2(prog_data[0]), .B1(\mem[189][0] ), .B2(n7418), 
        .Z(n1629) );
  NR2D0 U6410 ( .A1(n7570), .A2(n7422), .ZN(n7420) );
  INVD0 U6411 ( .I(n7420), .ZN(n7421) );
  OA22D0 U6412 ( .A1(n7421), .A2(prog_data[15]), .B1(\mem[190][15] ), .B2(
        n7420), .Z(n1628) );
  OA22D0 U6413 ( .A1(n7421), .A2(prog_data[14]), .B1(\mem[190][14] ), .B2(
        n7420), .Z(n1627) );
  OA22D0 U6414 ( .A1(n7421), .A2(prog_data[13]), .B1(\mem[190][13] ), .B2(
        n7420), .Z(n1626) );
  OA22D0 U6415 ( .A1(n7421), .A2(prog_data[12]), .B1(\mem[190][12] ), .B2(
        n7420), .Z(n1625) );
  OA22D0 U6416 ( .A1(n7421), .A2(prog_data[11]), .B1(\mem[190][11] ), .B2(
        n7420), .Z(n1624) );
  OA22D0 U6417 ( .A1(n7421), .A2(prog_data[10]), .B1(\mem[190][10] ), .B2(
        n7420), .Z(n1623) );
  OA22D0 U6418 ( .A1(n7421), .A2(prog_data[9]), .B1(\mem[190][9] ), .B2(n7420), 
        .Z(n1622) );
  OA22D0 U6419 ( .A1(n7421), .A2(prog_data[8]), .B1(\mem[190][8] ), .B2(n7420), 
        .Z(n1621) );
  OA22D0 U6420 ( .A1(n7421), .A2(prog_data[7]), .B1(\mem[190][7] ), .B2(n7420), 
        .Z(n1620) );
  OA22D0 U6421 ( .A1(n7421), .A2(prog_data[6]), .B1(\mem[190][6] ), .B2(n7420), 
        .Z(n1619) );
  OA22D0 U6422 ( .A1(n7421), .A2(prog_data[5]), .B1(\mem[190][5] ), .B2(n7420), 
        .Z(n1618) );
  OA22D0 U6423 ( .A1(n7421), .A2(prog_data[4]), .B1(\mem[190][4] ), .B2(n7420), 
        .Z(n1617) );
  OA22D0 U6424 ( .A1(n7421), .A2(prog_data[3]), .B1(\mem[190][3] ), .B2(n7420), 
        .Z(n1616) );
  OA22D0 U6425 ( .A1(n7421), .A2(prog_data[2]), .B1(\mem[190][2] ), .B2(n7420), 
        .Z(n1615) );
  OA22D0 U6426 ( .A1(n7421), .A2(prog_data[1]), .B1(\mem[190][1] ), .B2(n7420), 
        .Z(n1614) );
  OA22D0 U6427 ( .A1(n7421), .A2(prog_data[0]), .B1(\mem[190][0] ), .B2(n7420), 
        .Z(n1613) );
  NR2D0 U6428 ( .A1(n7574), .A2(n7422), .ZN(n7423) );
  INVD0 U6429 ( .I(n7423), .ZN(n7424) );
  OA22D0 U6430 ( .A1(n7424), .A2(prog_data[15]), .B1(\mem[191][15] ), .B2(
        n7423), .Z(n1612) );
  OA22D0 U6431 ( .A1(n7424), .A2(prog_data[14]), .B1(\mem[191][14] ), .B2(
        n7423), .Z(n1611) );
  OA22D0 U6432 ( .A1(n7424), .A2(prog_data[13]), .B1(\mem[191][13] ), .B2(
        n7423), .Z(n1610) );
  OA22D0 U6433 ( .A1(n7424), .A2(prog_data[12]), .B1(\mem[191][12] ), .B2(
        n7423), .Z(n1609) );
  OA22D0 U6434 ( .A1(n7424), .A2(prog_data[11]), .B1(\mem[191][11] ), .B2(
        n7423), .Z(n1608) );
  OA22D0 U6435 ( .A1(n7424), .A2(prog_data[10]), .B1(\mem[191][10] ), .B2(
        n7423), .Z(n1607) );
  OA22D0 U6436 ( .A1(n7424), .A2(prog_data[9]), .B1(\mem[191][9] ), .B2(n7423), 
        .Z(n1606) );
  OA22D0 U6437 ( .A1(n7424), .A2(prog_data[8]), .B1(\mem[191][8] ), .B2(n7423), 
        .Z(n1605) );
  OA22D0 U6438 ( .A1(n7424), .A2(prog_data[7]), .B1(\mem[191][7] ), .B2(n7423), 
        .Z(n1604) );
  OA22D0 U6439 ( .A1(n7424), .A2(prog_data[6]), .B1(\mem[191][6] ), .B2(n7423), 
        .Z(n1603) );
  OA22D0 U6440 ( .A1(n7424), .A2(prog_data[5]), .B1(\mem[191][5] ), .B2(n7423), 
        .Z(n1602) );
  OA22D0 U6441 ( .A1(n7424), .A2(prog_data[4]), .B1(\mem[191][4] ), .B2(n7423), 
        .Z(n1601) );
  OA22D0 U6442 ( .A1(n7424), .A2(prog_data[3]), .B1(\mem[191][3] ), .B2(n7423), 
        .Z(n1600) );
  OA22D0 U6443 ( .A1(n7424), .A2(prog_data[2]), .B1(\mem[191][2] ), .B2(n7423), 
        .Z(n1599) );
  OA22D0 U6444 ( .A1(n7424), .A2(prog_data[1]), .B1(\mem[191][1] ), .B2(n7423), 
        .Z(n1598) );
  OA22D0 U6445 ( .A1(n7424), .A2(prog_data[0]), .B1(\mem[191][0] ), .B2(n7423), 
        .Z(n1597) );
  IND3D0 U6446 ( .A1(n7458), .B1(prog_addr[6]), .B2(n7492), .ZN(n7455) );
  NR2D0 U6447 ( .A1(n7528), .A2(n7455), .ZN(n7425) );
  INVD0 U6448 ( .I(n7425), .ZN(n7426) );
  OA22D0 U6449 ( .A1(n7426), .A2(prog_data[15]), .B1(\mem[192][15] ), .B2(
        n7425), .Z(n1596) );
  OA22D0 U6450 ( .A1(n7426), .A2(prog_data[14]), .B1(\mem[192][14] ), .B2(
        n7425), .Z(n1595) );
  OA22D0 U6451 ( .A1(n7426), .A2(prog_data[13]), .B1(\mem[192][13] ), .B2(
        n7425), .Z(n1594) );
  OA22D0 U6452 ( .A1(n7426), .A2(prog_data[12]), .B1(\mem[192][12] ), .B2(
        n7425), .Z(n1593) );
  OA22D0 U6453 ( .A1(n7426), .A2(prog_data[11]), .B1(\mem[192][11] ), .B2(
        n7425), .Z(n1592) );
  OA22D0 U6454 ( .A1(n7426), .A2(prog_data[10]), .B1(\mem[192][10] ), .B2(
        n7425), .Z(n1591) );
  OA22D0 U6455 ( .A1(n7426), .A2(prog_data[9]), .B1(\mem[192][9] ), .B2(n7425), 
        .Z(n1590) );
  OA22D0 U6456 ( .A1(n7426), .A2(prog_data[8]), .B1(\mem[192][8] ), .B2(n7425), 
        .Z(n1589) );
  OA22D0 U6457 ( .A1(n7426), .A2(prog_data[7]), .B1(\mem[192][7] ), .B2(n7425), 
        .Z(n1588) );
  OA22D0 U6458 ( .A1(n7426), .A2(prog_data[6]), .B1(\mem[192][6] ), .B2(n7425), 
        .Z(n1587) );
  OA22D0 U6459 ( .A1(n7426), .A2(prog_data[5]), .B1(\mem[192][5] ), .B2(n7425), 
        .Z(n1586) );
  OA22D0 U6460 ( .A1(n7426), .A2(prog_data[4]), .B1(\mem[192][4] ), .B2(n7425), 
        .Z(n1585) );
  OA22D0 U6461 ( .A1(n7426), .A2(prog_data[3]), .B1(\mem[192][3] ), .B2(n7425), 
        .Z(n1584) );
  OA22D0 U6462 ( .A1(n7426), .A2(prog_data[2]), .B1(\mem[192][2] ), .B2(n7425), 
        .Z(n1583) );
  OA22D0 U6463 ( .A1(n7426), .A2(prog_data[1]), .B1(\mem[192][1] ), .B2(n7425), 
        .Z(n1582) );
  OA22D0 U6464 ( .A1(n7426), .A2(prog_data[0]), .B1(\mem[192][0] ), .B2(n7425), 
        .Z(n1581) );
  NR2D0 U6465 ( .A1(n7531), .A2(n7455), .ZN(n7427) );
  INVD0 U6466 ( .I(n7427), .ZN(n7428) );
  OA22D0 U6467 ( .A1(n7428), .A2(prog_data[15]), .B1(\mem[193][15] ), .B2(
        n7427), .Z(n1580) );
  OA22D0 U6468 ( .A1(n7428), .A2(prog_data[14]), .B1(\mem[193][14] ), .B2(
        n7427), .Z(n1579) );
  OA22D0 U6469 ( .A1(n7428), .A2(prog_data[13]), .B1(\mem[193][13] ), .B2(
        n7427), .Z(n1578) );
  OA22D0 U6470 ( .A1(n7428), .A2(prog_data[12]), .B1(\mem[193][12] ), .B2(
        n7427), .Z(n1577) );
  OA22D0 U6471 ( .A1(n7428), .A2(prog_data[11]), .B1(\mem[193][11] ), .B2(
        n7427), .Z(n1576) );
  OA22D0 U6472 ( .A1(n7428), .A2(prog_data[10]), .B1(\mem[193][10] ), .B2(
        n7427), .Z(n1575) );
  OA22D0 U6473 ( .A1(n7428), .A2(prog_data[9]), .B1(\mem[193][9] ), .B2(n7427), 
        .Z(n1574) );
  OA22D0 U6474 ( .A1(n7428), .A2(prog_data[8]), .B1(\mem[193][8] ), .B2(n7427), 
        .Z(n1573) );
  OA22D0 U6475 ( .A1(n7428), .A2(prog_data[7]), .B1(\mem[193][7] ), .B2(n7427), 
        .Z(n1572) );
  OA22D0 U6476 ( .A1(n7428), .A2(prog_data[6]), .B1(\mem[193][6] ), .B2(n7427), 
        .Z(n1571) );
  OA22D0 U6477 ( .A1(n7428), .A2(prog_data[5]), .B1(\mem[193][5] ), .B2(n7427), 
        .Z(n1570) );
  OA22D0 U6478 ( .A1(n7428), .A2(prog_data[4]), .B1(\mem[193][4] ), .B2(n7427), 
        .Z(n1569) );
  OA22D0 U6479 ( .A1(n7428), .A2(prog_data[3]), .B1(\mem[193][3] ), .B2(n7427), 
        .Z(n1568) );
  OA22D0 U6480 ( .A1(n7428), .A2(prog_data[2]), .B1(\mem[193][2] ), .B2(n7427), 
        .Z(n1567) );
  OA22D0 U6481 ( .A1(n7428), .A2(prog_data[1]), .B1(\mem[193][1] ), .B2(n7427), 
        .Z(n1566) );
  OA22D0 U6482 ( .A1(n7428), .A2(prog_data[0]), .B1(\mem[193][0] ), .B2(n7427), 
        .Z(n1565) );
  NR2D0 U6483 ( .A1(n7534), .A2(n7455), .ZN(n7429) );
  INVD0 U6484 ( .I(n7429), .ZN(n7430) );
  OA22D0 U6485 ( .A1(n7430), .A2(prog_data[15]), .B1(\mem[194][15] ), .B2(
        n7429), .Z(n1564) );
  OA22D0 U6486 ( .A1(n7430), .A2(prog_data[14]), .B1(\mem[194][14] ), .B2(
        n7429), .Z(n1563) );
  OA22D0 U6487 ( .A1(n7430), .A2(prog_data[13]), .B1(\mem[194][13] ), .B2(
        n7429), .Z(n1562) );
  OA22D0 U6488 ( .A1(n7430), .A2(prog_data[12]), .B1(\mem[194][12] ), .B2(
        n7429), .Z(n1561) );
  OA22D0 U6489 ( .A1(n7430), .A2(prog_data[11]), .B1(\mem[194][11] ), .B2(
        n7429), .Z(n1560) );
  OA22D0 U6490 ( .A1(n7430), .A2(prog_data[10]), .B1(\mem[194][10] ), .B2(
        n7429), .Z(n1559) );
  OA22D0 U6491 ( .A1(n7430), .A2(prog_data[9]), .B1(\mem[194][9] ), .B2(n7429), 
        .Z(n1558) );
  OA22D0 U6492 ( .A1(n7430), .A2(prog_data[8]), .B1(\mem[194][8] ), .B2(n7429), 
        .Z(n1557) );
  OA22D0 U6493 ( .A1(n7430), .A2(prog_data[7]), .B1(\mem[194][7] ), .B2(n7429), 
        .Z(n1556) );
  OA22D0 U6494 ( .A1(n7430), .A2(prog_data[6]), .B1(\mem[194][6] ), .B2(n7429), 
        .Z(n1555) );
  OA22D0 U6495 ( .A1(n7430), .A2(prog_data[5]), .B1(\mem[194][5] ), .B2(n7429), 
        .Z(n1554) );
  OA22D0 U6496 ( .A1(n7430), .A2(prog_data[4]), .B1(\mem[194][4] ), .B2(n7429), 
        .Z(n1553) );
  OA22D0 U6497 ( .A1(n7430), .A2(prog_data[3]), .B1(\mem[194][3] ), .B2(n7429), 
        .Z(n1552) );
  OA22D0 U6498 ( .A1(n7430), .A2(prog_data[2]), .B1(\mem[194][2] ), .B2(n7429), 
        .Z(n1551) );
  OA22D0 U6499 ( .A1(n7430), .A2(prog_data[1]), .B1(\mem[194][1] ), .B2(n7429), 
        .Z(n1550) );
  OA22D0 U6500 ( .A1(n7430), .A2(prog_data[0]), .B1(\mem[194][0] ), .B2(n7429), 
        .Z(n1549) );
  NR2D0 U6501 ( .A1(n7537), .A2(n7455), .ZN(n7431) );
  INVD0 U6502 ( .I(n7431), .ZN(n7432) );
  OA22D0 U6503 ( .A1(n7432), .A2(prog_data[15]), .B1(\mem[195][15] ), .B2(
        n7431), .Z(n1548) );
  OA22D0 U6504 ( .A1(n7432), .A2(prog_data[14]), .B1(\mem[195][14] ), .B2(
        n7431), .Z(n1547) );
  OA22D0 U6505 ( .A1(n7432), .A2(prog_data[13]), .B1(\mem[195][13] ), .B2(
        n7431), .Z(n1546) );
  OA22D0 U6506 ( .A1(n7432), .A2(prog_data[12]), .B1(\mem[195][12] ), .B2(
        n7431), .Z(n1545) );
  OA22D0 U6507 ( .A1(n7432), .A2(prog_data[11]), .B1(\mem[195][11] ), .B2(
        n7431), .Z(n1544) );
  OA22D0 U6508 ( .A1(n7432), .A2(prog_data[10]), .B1(\mem[195][10] ), .B2(
        n7431), .Z(n1543) );
  OA22D0 U6509 ( .A1(n7432), .A2(prog_data[9]), .B1(\mem[195][9] ), .B2(n7431), 
        .Z(n1542) );
  OA22D0 U6510 ( .A1(n7432), .A2(prog_data[8]), .B1(\mem[195][8] ), .B2(n7431), 
        .Z(n1541) );
  OA22D0 U6511 ( .A1(n7432), .A2(prog_data[7]), .B1(\mem[195][7] ), .B2(n7431), 
        .Z(n1540) );
  OA22D0 U6512 ( .A1(n7432), .A2(prog_data[6]), .B1(\mem[195][6] ), .B2(n7431), 
        .Z(n1539) );
  OA22D0 U6513 ( .A1(n7432), .A2(prog_data[5]), .B1(\mem[195][5] ), .B2(n7431), 
        .Z(n1538) );
  OA22D0 U6514 ( .A1(n7432), .A2(prog_data[4]), .B1(\mem[195][4] ), .B2(n7431), 
        .Z(n1537) );
  OA22D0 U6515 ( .A1(n7432), .A2(prog_data[3]), .B1(\mem[195][3] ), .B2(n7431), 
        .Z(n1536) );
  OA22D0 U6516 ( .A1(n7432), .A2(prog_data[2]), .B1(\mem[195][2] ), .B2(n7431), 
        .Z(n1535) );
  OA22D0 U6517 ( .A1(n7432), .A2(prog_data[1]), .B1(\mem[195][1] ), .B2(n7431), 
        .Z(n1534) );
  OA22D0 U6518 ( .A1(n7432), .A2(prog_data[0]), .B1(\mem[195][0] ), .B2(n7431), 
        .Z(n1533) );
  INVD0 U6519 ( .I(n7433), .ZN(n7434) );
  OA22D0 U6520 ( .A1(n7434), .A2(prog_data[15]), .B1(\mem[196][15] ), .B2(
        n7433), .Z(n1532) );
  OA22D0 U6521 ( .A1(n7434), .A2(prog_data[14]), .B1(\mem[196][14] ), .B2(
        n7433), .Z(n1531) );
  OA22D0 U6522 ( .A1(n7434), .A2(prog_data[13]), .B1(\mem[196][13] ), .B2(
        n7433), .Z(n1530) );
  OA22D0 U6523 ( .A1(n7434), .A2(prog_data[12]), .B1(\mem[196][12] ), .B2(
        n7433), .Z(n1529) );
  OA22D0 U6524 ( .A1(n7434), .A2(prog_data[11]), .B1(\mem[196][11] ), .B2(
        n7433), .Z(n1528) );
  OA22D0 U6525 ( .A1(n7434), .A2(prog_data[10]), .B1(\mem[196][10] ), .B2(
        n7433), .Z(n1527) );
  OA22D0 U6526 ( .A1(n7434), .A2(prog_data[9]), .B1(\mem[196][9] ), .B2(n7433), 
        .Z(n1526) );
  OA22D0 U6527 ( .A1(n7434), .A2(prog_data[8]), .B1(\mem[196][8] ), .B2(n7433), 
        .Z(n1525) );
  OA22D0 U6528 ( .A1(n7434), .A2(prog_data[7]), .B1(\mem[196][7] ), .B2(n7433), 
        .Z(n1524) );
  OA22D0 U6529 ( .A1(n7434), .A2(prog_data[6]), .B1(\mem[196][6] ), .B2(n7433), 
        .Z(n1523) );
  OA22D0 U6530 ( .A1(n7434), .A2(prog_data[5]), .B1(\mem[196][5] ), .B2(n7433), 
        .Z(n1522) );
  OA22D0 U6531 ( .A1(n7434), .A2(prog_data[4]), .B1(\mem[196][4] ), .B2(n7433), 
        .Z(n1521) );
  OA22D0 U6532 ( .A1(n7434), .A2(prog_data[3]), .B1(\mem[196][3] ), .B2(n7433), 
        .Z(n1520) );
  OA22D0 U6533 ( .A1(n7434), .A2(prog_data[2]), .B1(\mem[196][2] ), .B2(n7433), 
        .Z(n1519) );
  OA22D0 U6534 ( .A1(n7434), .A2(prog_data[1]), .B1(\mem[196][1] ), .B2(n7433), 
        .Z(n1518) );
  OA22D0 U6535 ( .A1(n7434), .A2(prog_data[0]), .B1(\mem[196][0] ), .B2(n7433), 
        .Z(n1517) );
  NR2D0 U6536 ( .A1(n7543), .A2(n7455), .ZN(n7435) );
  INVD0 U6537 ( .I(n7435), .ZN(n7436) );
  OA22D0 U6538 ( .A1(n7436), .A2(prog_data[15]), .B1(\mem[197][15] ), .B2(
        n7435), .Z(n1516) );
  OA22D0 U6539 ( .A1(n7436), .A2(prog_data[14]), .B1(\mem[197][14] ), .B2(
        n7435), .Z(n1515) );
  OA22D0 U6540 ( .A1(n7436), .A2(prog_data[13]), .B1(\mem[197][13] ), .B2(
        n7435), .Z(n1514) );
  OA22D0 U6541 ( .A1(n7436), .A2(prog_data[12]), .B1(\mem[197][12] ), .B2(
        n7435), .Z(n1513) );
  OA22D0 U6542 ( .A1(n7436), .A2(prog_data[11]), .B1(\mem[197][11] ), .B2(
        n7435), .Z(n1512) );
  OA22D0 U6543 ( .A1(n7436), .A2(prog_data[10]), .B1(\mem[197][10] ), .B2(
        n7435), .Z(n1511) );
  OA22D0 U6544 ( .A1(n7436), .A2(prog_data[9]), .B1(\mem[197][9] ), .B2(n7435), 
        .Z(n1510) );
  OA22D0 U6545 ( .A1(n7436), .A2(prog_data[8]), .B1(\mem[197][8] ), .B2(n7435), 
        .Z(n1509) );
  OA22D0 U6546 ( .A1(n7436), .A2(prog_data[7]), .B1(\mem[197][7] ), .B2(n7435), 
        .Z(n1508) );
  OA22D0 U6547 ( .A1(n7436), .A2(prog_data[6]), .B1(\mem[197][6] ), .B2(n7435), 
        .Z(n1507) );
  OA22D0 U6548 ( .A1(n7436), .A2(prog_data[5]), .B1(\mem[197][5] ), .B2(n7435), 
        .Z(n1506) );
  OA22D0 U6549 ( .A1(n7436), .A2(prog_data[4]), .B1(\mem[197][4] ), .B2(n7435), 
        .Z(n1505) );
  OA22D0 U6550 ( .A1(n7436), .A2(prog_data[3]), .B1(\mem[197][3] ), .B2(n7435), 
        .Z(n1504) );
  OA22D0 U6551 ( .A1(n7436), .A2(prog_data[2]), .B1(\mem[197][2] ), .B2(n7435), 
        .Z(n1503) );
  OA22D0 U6552 ( .A1(n7436), .A2(prog_data[1]), .B1(\mem[197][1] ), .B2(n7435), 
        .Z(n1502) );
  OA22D0 U6553 ( .A1(n7436), .A2(prog_data[0]), .B1(\mem[197][0] ), .B2(n7435), 
        .Z(n1501) );
  NR2D0 U6554 ( .A1(n7546), .A2(n7455), .ZN(n7437) );
  INVD0 U6555 ( .I(n7437), .ZN(n7438) );
  OA22D0 U6556 ( .A1(n7438), .A2(prog_data[15]), .B1(\mem[198][15] ), .B2(
        n7437), .Z(n1500) );
  OA22D0 U6557 ( .A1(n7438), .A2(prog_data[14]), .B1(\mem[198][14] ), .B2(
        n7437), .Z(n1499) );
  OA22D0 U6558 ( .A1(n7438), .A2(prog_data[13]), .B1(\mem[198][13] ), .B2(
        n7437), .Z(n1498) );
  OA22D0 U6559 ( .A1(n7438), .A2(prog_data[12]), .B1(\mem[198][12] ), .B2(
        n7437), .Z(n1497) );
  OA22D0 U6560 ( .A1(n7438), .A2(prog_data[11]), .B1(\mem[198][11] ), .B2(
        n7437), .Z(n1496) );
  OA22D0 U6561 ( .A1(n7438), .A2(prog_data[10]), .B1(\mem[198][10] ), .B2(
        n7437), .Z(n1495) );
  OA22D0 U6562 ( .A1(n7438), .A2(prog_data[9]), .B1(\mem[198][9] ), .B2(n7437), 
        .Z(n1494) );
  OA22D0 U6563 ( .A1(n7438), .A2(prog_data[8]), .B1(\mem[198][8] ), .B2(n7437), 
        .Z(n1493) );
  OA22D0 U6564 ( .A1(n7438), .A2(prog_data[7]), .B1(\mem[198][7] ), .B2(n7437), 
        .Z(n1492) );
  OA22D0 U6565 ( .A1(n7438), .A2(prog_data[6]), .B1(\mem[198][6] ), .B2(n7437), 
        .Z(n1491) );
  OA22D0 U6566 ( .A1(n7438), .A2(prog_data[5]), .B1(\mem[198][5] ), .B2(n7437), 
        .Z(n1490) );
  OA22D0 U6567 ( .A1(n7438), .A2(prog_data[4]), .B1(\mem[198][4] ), .B2(n7437), 
        .Z(n1489) );
  OA22D0 U6568 ( .A1(n7438), .A2(prog_data[3]), .B1(\mem[198][3] ), .B2(n7437), 
        .Z(n1488) );
  OA22D0 U6569 ( .A1(n7438), .A2(prog_data[2]), .B1(\mem[198][2] ), .B2(n7437), 
        .Z(n1487) );
  OA22D0 U6570 ( .A1(n7438), .A2(prog_data[1]), .B1(\mem[198][1] ), .B2(n7437), 
        .Z(n1486) );
  OA22D0 U6571 ( .A1(n7438), .A2(prog_data[0]), .B1(\mem[198][0] ), .B2(n7437), 
        .Z(n1485) );
  NR2D0 U6572 ( .A1(n7549), .A2(n7455), .ZN(n7439) );
  INVD0 U6573 ( .I(n7439), .ZN(n7440) );
  OA22D0 U6574 ( .A1(n7440), .A2(prog_data[15]), .B1(\mem[199][15] ), .B2(
        n7439), .Z(n1484) );
  OA22D0 U6575 ( .A1(n7440), .A2(prog_data[14]), .B1(\mem[199][14] ), .B2(
        n7439), .Z(n1483) );
  OA22D0 U6576 ( .A1(n7440), .A2(prog_data[13]), .B1(\mem[199][13] ), .B2(
        n7439), .Z(n1482) );
  OA22D0 U6577 ( .A1(n7440), .A2(prog_data[12]), .B1(\mem[199][12] ), .B2(
        n7439), .Z(n1481) );
  OA22D0 U6578 ( .A1(n7440), .A2(prog_data[11]), .B1(\mem[199][11] ), .B2(
        n7439), .Z(n1480) );
  OA22D0 U6579 ( .A1(n7440), .A2(prog_data[10]), .B1(\mem[199][10] ), .B2(
        n7439), .Z(n1479) );
  OA22D0 U6580 ( .A1(n7440), .A2(prog_data[9]), .B1(\mem[199][9] ), .B2(n7439), 
        .Z(n1478) );
  OA22D0 U6581 ( .A1(n7440), .A2(prog_data[8]), .B1(\mem[199][8] ), .B2(n7439), 
        .Z(n1477) );
  OA22D0 U6582 ( .A1(n7440), .A2(prog_data[7]), .B1(\mem[199][7] ), .B2(n7439), 
        .Z(n1476) );
  OA22D0 U6583 ( .A1(n7440), .A2(prog_data[6]), .B1(\mem[199][6] ), .B2(n7439), 
        .Z(n1475) );
  OA22D0 U6584 ( .A1(n7440), .A2(prog_data[5]), .B1(\mem[199][5] ), .B2(n7439), 
        .Z(n1474) );
  OA22D0 U6585 ( .A1(n7440), .A2(prog_data[4]), .B1(\mem[199][4] ), .B2(n7439), 
        .Z(n1473) );
  OA22D0 U6586 ( .A1(n7440), .A2(prog_data[3]), .B1(\mem[199][3] ), .B2(n7439), 
        .Z(n1472) );
  OA22D0 U6587 ( .A1(n7440), .A2(prog_data[2]), .B1(\mem[199][2] ), .B2(n7439), 
        .Z(n1471) );
  OA22D0 U6588 ( .A1(n7440), .A2(prog_data[1]), .B1(\mem[199][1] ), .B2(n7439), 
        .Z(n1470) );
  OA22D0 U6589 ( .A1(n7440), .A2(prog_data[0]), .B1(\mem[199][0] ), .B2(n7439), 
        .Z(n1469) );
  NR2D0 U6590 ( .A1(n7552), .A2(n7455), .ZN(n7441) );
  INVD0 U6591 ( .I(n7441), .ZN(n7442) );
  OA22D0 U6592 ( .A1(n7442), .A2(prog_data[15]), .B1(\mem[200][15] ), .B2(
        n7441), .Z(n1468) );
  OA22D0 U6593 ( .A1(n7442), .A2(prog_data[14]), .B1(\mem[200][14] ), .B2(
        n7441), .Z(n1467) );
  OA22D0 U6594 ( .A1(n7442), .A2(prog_data[13]), .B1(\mem[200][13] ), .B2(
        n7441), .Z(n1466) );
  OA22D0 U6595 ( .A1(n7442), .A2(prog_data[12]), .B1(\mem[200][12] ), .B2(
        n7441), .Z(n1465) );
  OA22D0 U6596 ( .A1(n7442), .A2(prog_data[11]), .B1(\mem[200][11] ), .B2(
        n7441), .Z(n1464) );
  OA22D0 U6597 ( .A1(n7442), .A2(prog_data[10]), .B1(\mem[200][10] ), .B2(
        n7441), .Z(n1463) );
  OA22D0 U6598 ( .A1(n7442), .A2(prog_data[9]), .B1(\mem[200][9] ), .B2(n7441), 
        .Z(n1462) );
  OA22D0 U6599 ( .A1(n7442), .A2(prog_data[8]), .B1(\mem[200][8] ), .B2(n7441), 
        .Z(n1461) );
  OA22D0 U6600 ( .A1(n7442), .A2(prog_data[7]), .B1(\mem[200][7] ), .B2(n7441), 
        .Z(n1460) );
  OA22D0 U6601 ( .A1(n7442), .A2(prog_data[6]), .B1(\mem[200][6] ), .B2(n7441), 
        .Z(n1459) );
  OA22D0 U6602 ( .A1(n7442), .A2(prog_data[5]), .B1(\mem[200][5] ), .B2(n7441), 
        .Z(n1458) );
  OA22D0 U6603 ( .A1(n7442), .A2(prog_data[4]), .B1(\mem[200][4] ), .B2(n7441), 
        .Z(n1457) );
  OA22D0 U6604 ( .A1(n7442), .A2(prog_data[3]), .B1(\mem[200][3] ), .B2(n7441), 
        .Z(n1456) );
  OA22D0 U6605 ( .A1(n7442), .A2(prog_data[2]), .B1(\mem[200][2] ), .B2(n7441), 
        .Z(n1455) );
  OA22D0 U6606 ( .A1(n7442), .A2(prog_data[1]), .B1(\mem[200][1] ), .B2(n7441), 
        .Z(n1454) );
  OA22D0 U6607 ( .A1(n7442), .A2(prog_data[0]), .B1(\mem[200][0] ), .B2(n7441), 
        .Z(n1453) );
  NR2D0 U6608 ( .A1(n7555), .A2(n7455), .ZN(n7443) );
  INVD0 U6609 ( .I(n7443), .ZN(n7444) );
  OA22D0 U6610 ( .A1(n7444), .A2(prog_data[15]), .B1(\mem[201][15] ), .B2(
        n7443), .Z(n1452) );
  OA22D0 U6611 ( .A1(n7444), .A2(prog_data[14]), .B1(\mem[201][14] ), .B2(
        n7443), .Z(n1451) );
  OA22D0 U6612 ( .A1(n7444), .A2(prog_data[13]), .B1(\mem[201][13] ), .B2(
        n7443), .Z(n1450) );
  OA22D0 U6613 ( .A1(n7444), .A2(prog_data[12]), .B1(\mem[201][12] ), .B2(
        n7443), .Z(n1449) );
  OA22D0 U6614 ( .A1(n7444), .A2(prog_data[11]), .B1(\mem[201][11] ), .B2(
        n7443), .Z(n1448) );
  OA22D0 U6615 ( .A1(n7444), .A2(prog_data[10]), .B1(\mem[201][10] ), .B2(
        n7443), .Z(n1447) );
  OA22D0 U6616 ( .A1(n7444), .A2(prog_data[9]), .B1(\mem[201][9] ), .B2(n7443), 
        .Z(n1446) );
  OA22D0 U6617 ( .A1(n7444), .A2(prog_data[8]), .B1(\mem[201][8] ), .B2(n7443), 
        .Z(n1445) );
  OA22D0 U6618 ( .A1(n7444), .A2(prog_data[7]), .B1(\mem[201][7] ), .B2(n7443), 
        .Z(n1444) );
  OA22D0 U6619 ( .A1(n7444), .A2(prog_data[6]), .B1(\mem[201][6] ), .B2(n7443), 
        .Z(n1443) );
  OA22D0 U6620 ( .A1(n7444), .A2(prog_data[5]), .B1(\mem[201][5] ), .B2(n7443), 
        .Z(n1442) );
  OA22D0 U6621 ( .A1(n7444), .A2(prog_data[4]), .B1(\mem[201][4] ), .B2(n7443), 
        .Z(n1441) );
  OA22D0 U6622 ( .A1(n7444), .A2(prog_data[3]), .B1(\mem[201][3] ), .B2(n7443), 
        .Z(n1440) );
  OA22D0 U6623 ( .A1(n7444), .A2(prog_data[2]), .B1(\mem[201][2] ), .B2(n7443), 
        .Z(n1439) );
  OA22D0 U6624 ( .A1(n7444), .A2(prog_data[1]), .B1(\mem[201][1] ), .B2(n7443), 
        .Z(n1438) );
  OA22D0 U6625 ( .A1(n7444), .A2(prog_data[0]), .B1(\mem[201][0] ), .B2(n7443), 
        .Z(n1437) );
  NR2D0 U6626 ( .A1(n7558), .A2(n7455), .ZN(n7445) );
  INVD0 U6627 ( .I(n7445), .ZN(n7446) );
  OA22D0 U6628 ( .A1(n7446), .A2(prog_data[15]), .B1(\mem[202][15] ), .B2(
        n7445), .Z(n1436) );
  OA22D0 U6629 ( .A1(n7446), .A2(prog_data[14]), .B1(\mem[202][14] ), .B2(
        n7445), .Z(n1435) );
  OA22D0 U6630 ( .A1(n7446), .A2(prog_data[13]), .B1(\mem[202][13] ), .B2(
        n7445), .Z(n1434) );
  OA22D0 U6631 ( .A1(n7446), .A2(prog_data[12]), .B1(\mem[202][12] ), .B2(
        n7445), .Z(n1433) );
  OA22D0 U6632 ( .A1(n7446), .A2(prog_data[11]), .B1(\mem[202][11] ), .B2(
        n7445), .Z(n1432) );
  OA22D0 U6633 ( .A1(n7446), .A2(prog_data[10]), .B1(\mem[202][10] ), .B2(
        n7445), .Z(n1431) );
  OA22D0 U6634 ( .A1(n7446), .A2(prog_data[9]), .B1(\mem[202][9] ), .B2(n7445), 
        .Z(n1430) );
  OA22D0 U6635 ( .A1(n7446), .A2(prog_data[8]), .B1(\mem[202][8] ), .B2(n7445), 
        .Z(n1429) );
  OA22D0 U6636 ( .A1(n7446), .A2(prog_data[7]), .B1(\mem[202][7] ), .B2(n7445), 
        .Z(n1428) );
  OA22D0 U6637 ( .A1(n7446), .A2(prog_data[6]), .B1(\mem[202][6] ), .B2(n7445), 
        .Z(n1427) );
  OA22D0 U6638 ( .A1(n7446), .A2(prog_data[5]), .B1(\mem[202][5] ), .B2(n7445), 
        .Z(n1426) );
  OA22D0 U6639 ( .A1(n7446), .A2(prog_data[4]), .B1(\mem[202][4] ), .B2(n7445), 
        .Z(n1425) );
  OA22D0 U6640 ( .A1(n7446), .A2(prog_data[3]), .B1(\mem[202][3] ), .B2(n7445), 
        .Z(n1424) );
  OA22D0 U6641 ( .A1(n7446), .A2(prog_data[2]), .B1(\mem[202][2] ), .B2(n7445), 
        .Z(n1423) );
  OA22D0 U6642 ( .A1(n7446), .A2(prog_data[1]), .B1(\mem[202][1] ), .B2(n7445), 
        .Z(n1422) );
  OA22D0 U6643 ( .A1(n7446), .A2(prog_data[0]), .B1(\mem[202][0] ), .B2(n7445), 
        .Z(n1421) );
  NR2D0 U6644 ( .A1(n7561), .A2(n7455), .ZN(n7447) );
  INVD0 U6645 ( .I(n7447), .ZN(n7448) );
  OA22D0 U6646 ( .A1(n7448), .A2(prog_data[15]), .B1(\mem[203][15] ), .B2(
        n7447), .Z(n1420) );
  OA22D0 U6647 ( .A1(n7448), .A2(prog_data[14]), .B1(\mem[203][14] ), .B2(
        n7447), .Z(n1419) );
  OA22D0 U6648 ( .A1(n7448), .A2(prog_data[13]), .B1(\mem[203][13] ), .B2(
        n7447), .Z(n1418) );
  OA22D0 U6649 ( .A1(n7448), .A2(prog_data[12]), .B1(\mem[203][12] ), .B2(
        n7447), .Z(n1417) );
  OA22D0 U6650 ( .A1(n7448), .A2(prog_data[11]), .B1(\mem[203][11] ), .B2(
        n7447), .Z(n1416) );
  OA22D0 U6651 ( .A1(n7448), .A2(prog_data[10]), .B1(\mem[203][10] ), .B2(
        n7447), .Z(n1415) );
  OA22D0 U6652 ( .A1(n7448), .A2(prog_data[9]), .B1(\mem[203][9] ), .B2(n7447), 
        .Z(n1414) );
  OA22D0 U6653 ( .A1(n7448), .A2(prog_data[8]), .B1(\mem[203][8] ), .B2(n7447), 
        .Z(n1413) );
  OA22D0 U6654 ( .A1(n7448), .A2(prog_data[7]), .B1(\mem[203][7] ), .B2(n7447), 
        .Z(n1412) );
  OA22D0 U6655 ( .A1(n7448), .A2(prog_data[6]), .B1(\mem[203][6] ), .B2(n7447), 
        .Z(n1411) );
  OA22D0 U6656 ( .A1(n7448), .A2(prog_data[5]), .B1(\mem[203][5] ), .B2(n7447), 
        .Z(n1410) );
  OA22D0 U6657 ( .A1(n7448), .A2(prog_data[4]), .B1(\mem[203][4] ), .B2(n7447), 
        .Z(n1409) );
  OA22D0 U6658 ( .A1(n7448), .A2(prog_data[3]), .B1(\mem[203][3] ), .B2(n7447), 
        .Z(n1408) );
  OA22D0 U6659 ( .A1(n7448), .A2(prog_data[2]), .B1(\mem[203][2] ), .B2(n7447), 
        .Z(n1407) );
  OA22D0 U6660 ( .A1(n7448), .A2(prog_data[1]), .B1(\mem[203][1] ), .B2(n7447), 
        .Z(n1406) );
  OA22D0 U6661 ( .A1(n7448), .A2(prog_data[0]), .B1(\mem[203][0] ), .B2(n7447), 
        .Z(n1405) );
  NR2D0 U6662 ( .A1(n7564), .A2(n7455), .ZN(n7449) );
  OA22D0 U6663 ( .A1(n7450), .A2(prog_data[15]), .B1(\mem[204][15] ), .B2(
        n7449), .Z(n1404) );
  OA22D0 U6664 ( .A1(n7450), .A2(prog_data[14]), .B1(\mem[204][14] ), .B2(
        n7449), .Z(n1403) );
  OA22D0 U6665 ( .A1(n7450), .A2(prog_data[13]), .B1(\mem[204][13] ), .B2(
        n7449), .Z(n1402) );
  OA22D0 U6666 ( .A1(n7450), .A2(prog_data[12]), .B1(\mem[204][12] ), .B2(
        n7449), .Z(n1401) );
  OA22D0 U6667 ( .A1(n7450), .A2(prog_data[11]), .B1(\mem[204][11] ), .B2(
        n7449), .Z(n1400) );
  OA22D0 U6668 ( .A1(n7450), .A2(prog_data[10]), .B1(\mem[204][10] ), .B2(
        n7449), .Z(n1399) );
  OA22D0 U6669 ( .A1(n7450), .A2(prog_data[9]), .B1(\mem[204][9] ), .B2(n7449), 
        .Z(n1398) );
  OA22D0 U6670 ( .A1(n7450), .A2(prog_data[8]), .B1(\mem[204][8] ), .B2(n7449), 
        .Z(n1397) );
  OA22D0 U6671 ( .A1(n7450), .A2(prog_data[7]), .B1(\mem[204][7] ), .B2(n7449), 
        .Z(n1396) );
  OA22D0 U6672 ( .A1(n7450), .A2(prog_data[6]), .B1(\mem[204][6] ), .B2(n7449), 
        .Z(n1395) );
  OA22D0 U6673 ( .A1(n7450), .A2(prog_data[5]), .B1(\mem[204][5] ), .B2(n7449), 
        .Z(n1394) );
  OA22D0 U6674 ( .A1(n7450), .A2(prog_data[4]), .B1(\mem[204][4] ), .B2(n7449), 
        .Z(n1393) );
  OA22D0 U6675 ( .A1(n7450), .A2(prog_data[3]), .B1(\mem[204][3] ), .B2(n7449), 
        .Z(n1392) );
  OA22D0 U6676 ( .A1(n7450), .A2(prog_data[2]), .B1(\mem[204][2] ), .B2(n7449), 
        .Z(n1391) );
  OA22D0 U6677 ( .A1(n7450), .A2(prog_data[1]), .B1(\mem[204][1] ), .B2(n7449), 
        .Z(n1390) );
  OA22D0 U6678 ( .A1(n7450), .A2(prog_data[0]), .B1(\mem[204][0] ), .B2(n7449), 
        .Z(n1389) );
  NR2D0 U6679 ( .A1(n7567), .A2(n7455), .ZN(n7451) );
  INVD0 U6680 ( .I(n7451), .ZN(n7452) );
  OA22D0 U6681 ( .A1(n7452), .A2(prog_data[15]), .B1(\mem[205][15] ), .B2(
        n7451), .Z(n1388) );
  OA22D0 U6682 ( .A1(n7452), .A2(prog_data[14]), .B1(\mem[205][14] ), .B2(
        n7451), .Z(n1387) );
  OA22D0 U6683 ( .A1(n7452), .A2(prog_data[13]), .B1(\mem[205][13] ), .B2(
        n7451), .Z(n1386) );
  OA22D0 U6684 ( .A1(n7452), .A2(prog_data[12]), .B1(\mem[205][12] ), .B2(
        n7451), .Z(n1385) );
  OA22D0 U6685 ( .A1(n7452), .A2(prog_data[11]), .B1(\mem[205][11] ), .B2(
        n7451), .Z(n1384) );
  OA22D0 U6686 ( .A1(n7452), .A2(prog_data[10]), .B1(\mem[205][10] ), .B2(
        n7451), .Z(n1383) );
  OA22D0 U6687 ( .A1(n7452), .A2(prog_data[9]), .B1(\mem[205][9] ), .B2(n7451), 
        .Z(n1382) );
  OA22D0 U6688 ( .A1(n7452), .A2(prog_data[8]), .B1(\mem[205][8] ), .B2(n7451), 
        .Z(n1381) );
  OA22D0 U6689 ( .A1(n7452), .A2(prog_data[7]), .B1(\mem[205][7] ), .B2(n7451), 
        .Z(n1380) );
  OA22D0 U6690 ( .A1(n7452), .A2(prog_data[6]), .B1(\mem[205][6] ), .B2(n7451), 
        .Z(n1379) );
  OA22D0 U6691 ( .A1(n7452), .A2(prog_data[5]), .B1(\mem[205][5] ), .B2(n7451), 
        .Z(n1378) );
  OA22D0 U6692 ( .A1(n7452), .A2(prog_data[4]), .B1(\mem[205][4] ), .B2(n7451), 
        .Z(n1377) );
  OA22D0 U6693 ( .A1(n7452), .A2(prog_data[3]), .B1(\mem[205][3] ), .B2(n7451), 
        .Z(n1376) );
  OA22D0 U6694 ( .A1(n7452), .A2(prog_data[2]), .B1(\mem[205][2] ), .B2(n7451), 
        .Z(n1375) );
  OA22D0 U6695 ( .A1(n7452), .A2(prog_data[1]), .B1(\mem[205][1] ), .B2(n7451), 
        .Z(n1374) );
  OA22D0 U6696 ( .A1(n7452), .A2(prog_data[0]), .B1(\mem[205][0] ), .B2(n7451), 
        .Z(n1373) );
  NR2D0 U6697 ( .A1(n7570), .A2(n7455), .ZN(n7453) );
  INVD0 U6698 ( .I(n7453), .ZN(n7454) );
  OA22D0 U6699 ( .A1(n7454), .A2(prog_data[15]), .B1(\mem[206][15] ), .B2(
        n7453), .Z(n1372) );
  OA22D0 U6700 ( .A1(n7454), .A2(prog_data[14]), .B1(\mem[206][14] ), .B2(
        n7453), .Z(n1371) );
  OA22D0 U6701 ( .A1(n7454), .A2(prog_data[13]), .B1(\mem[206][13] ), .B2(
        n7453), .Z(n1370) );
  OA22D0 U6702 ( .A1(n7454), .A2(prog_data[12]), .B1(\mem[206][12] ), .B2(
        n7453), .Z(n1369) );
  OA22D0 U6703 ( .A1(n7454), .A2(prog_data[11]), .B1(\mem[206][11] ), .B2(
        n7453), .Z(n1368) );
  OA22D0 U6704 ( .A1(n7454), .A2(prog_data[10]), .B1(\mem[206][10] ), .B2(
        n7453), .Z(n1367) );
  OA22D0 U6705 ( .A1(n7454), .A2(prog_data[9]), .B1(\mem[206][9] ), .B2(n7453), 
        .Z(n1366) );
  OA22D0 U6706 ( .A1(n7454), .A2(prog_data[8]), .B1(\mem[206][8] ), .B2(n7453), 
        .Z(n1365) );
  OA22D0 U6707 ( .A1(n7454), .A2(prog_data[7]), .B1(\mem[206][7] ), .B2(n7453), 
        .Z(n1364) );
  OA22D0 U6708 ( .A1(n7454), .A2(prog_data[6]), .B1(\mem[206][6] ), .B2(n7453), 
        .Z(n1363) );
  OA22D0 U6709 ( .A1(n7454), .A2(prog_data[5]), .B1(\mem[206][5] ), .B2(n7453), 
        .Z(n1362) );
  OA22D0 U6710 ( .A1(n7454), .A2(prog_data[4]), .B1(\mem[206][4] ), .B2(n7453), 
        .Z(n1361) );
  OA22D0 U6711 ( .A1(n7454), .A2(prog_data[3]), .B1(\mem[206][3] ), .B2(n7453), 
        .Z(n1360) );
  OA22D0 U6712 ( .A1(n7454), .A2(prog_data[2]), .B1(\mem[206][2] ), .B2(n7453), 
        .Z(n1359) );
  OA22D0 U6713 ( .A1(n7454), .A2(prog_data[1]), .B1(\mem[206][1] ), .B2(n7453), 
        .Z(n1358) );
  OA22D0 U6714 ( .A1(n7454), .A2(prog_data[0]), .B1(\mem[206][0] ), .B2(n7453), 
        .Z(n1357) );
  NR2D0 U6715 ( .A1(n7574), .A2(n7455), .ZN(n7456) );
  INVD0 U6716 ( .I(n7456), .ZN(n7457) );
  OA22D0 U6717 ( .A1(n7457), .A2(prog_data[15]), .B1(\mem[207][15] ), .B2(
        n7456), .Z(n1356) );
  OA22D0 U6718 ( .A1(n7457), .A2(prog_data[14]), .B1(\mem[207][14] ), .B2(
        n7456), .Z(n1355) );
  OA22D0 U6719 ( .A1(n7457), .A2(prog_data[13]), .B1(\mem[207][13] ), .B2(
        n7456), .Z(n1354) );
  OA22D0 U6720 ( .A1(n7457), .A2(prog_data[12]), .B1(\mem[207][12] ), .B2(
        n7456), .Z(n1353) );
  OA22D0 U6721 ( .A1(n7457), .A2(prog_data[11]), .B1(\mem[207][11] ), .B2(
        n7456), .Z(n1352) );
  OA22D0 U6722 ( .A1(n7457), .A2(prog_data[10]), .B1(\mem[207][10] ), .B2(
        n7456), .Z(n1351) );
  OA22D0 U6723 ( .A1(n7457), .A2(prog_data[9]), .B1(\mem[207][9] ), .B2(n7456), 
        .Z(n1350) );
  OA22D0 U6724 ( .A1(n7457), .A2(prog_data[8]), .B1(\mem[207][8] ), .B2(n7456), 
        .Z(n1349) );
  OA22D0 U6725 ( .A1(n7457), .A2(prog_data[7]), .B1(\mem[207][7] ), .B2(n7456), 
        .Z(n1348) );
  OA22D0 U6726 ( .A1(n7457), .A2(prog_data[6]), .B1(\mem[207][6] ), .B2(n7456), 
        .Z(n1347) );
  OA22D0 U6727 ( .A1(n7457), .A2(prog_data[5]), .B1(\mem[207][5] ), .B2(n7456), 
        .Z(n1346) );
  OA22D0 U6728 ( .A1(n7457), .A2(prog_data[4]), .B1(\mem[207][4] ), .B2(n7456), 
        .Z(n1345) );
  OA22D0 U6729 ( .A1(n7457), .A2(prog_data[3]), .B1(\mem[207][3] ), .B2(n7456), 
        .Z(n1344) );
  OA22D0 U6730 ( .A1(n7457), .A2(prog_data[2]), .B1(\mem[207][2] ), .B2(n7456), 
        .Z(n1343) );
  OA22D0 U6731 ( .A1(n7457), .A2(prog_data[1]), .B1(\mem[207][1] ), .B2(n7456), 
        .Z(n1342) );
  OA22D0 U6732 ( .A1(n7457), .A2(prog_data[0]), .B1(\mem[207][0] ), .B2(n7456), 
        .Z(n1341) );
  IND3D0 U6733 ( .A1(n7458), .B1(prog_addr[6]), .B2(n7526), .ZN(n7489) );
  NR2D0 U6734 ( .A1(n7528), .A2(n7489), .ZN(n7459) );
  INVD0 U6735 ( .I(n7459), .ZN(n7460) );
  OA22D0 U6736 ( .A1(n7460), .A2(prog_data[15]), .B1(\mem[208][15] ), .B2(
        n7459), .Z(n1340) );
  OA22D0 U6737 ( .A1(n7460), .A2(prog_data[14]), .B1(\mem[208][14] ), .B2(
        n7459), .Z(n1339) );
  OA22D0 U6738 ( .A1(n7460), .A2(prog_data[13]), .B1(\mem[208][13] ), .B2(
        n7459), .Z(n1338) );
  OA22D0 U6739 ( .A1(n7460), .A2(prog_data[12]), .B1(\mem[208][12] ), .B2(
        n7459), .Z(n1337) );
  OA22D0 U6740 ( .A1(n7460), .A2(prog_data[11]), .B1(\mem[208][11] ), .B2(
        n7459), .Z(n1336) );
  OA22D0 U6741 ( .A1(n7460), .A2(prog_data[10]), .B1(\mem[208][10] ), .B2(
        n7459), .Z(n1335) );
  OA22D0 U6742 ( .A1(n7460), .A2(prog_data[9]), .B1(\mem[208][9] ), .B2(n7459), 
        .Z(n1334) );
  OA22D0 U6743 ( .A1(n7460), .A2(prog_data[8]), .B1(\mem[208][8] ), .B2(n7459), 
        .Z(n1333) );
  OA22D0 U6744 ( .A1(n7460), .A2(prog_data[7]), .B1(\mem[208][7] ), .B2(n7459), 
        .Z(n1332) );
  OA22D0 U6745 ( .A1(n7460), .A2(prog_data[6]), .B1(\mem[208][6] ), .B2(n7459), 
        .Z(n1331) );
  OA22D0 U6746 ( .A1(n7460), .A2(prog_data[5]), .B1(\mem[208][5] ), .B2(n7459), 
        .Z(n1330) );
  OA22D0 U6747 ( .A1(n7460), .A2(prog_data[4]), .B1(\mem[208][4] ), .B2(n7459), 
        .Z(n1329) );
  OA22D0 U6748 ( .A1(n7460), .A2(prog_data[3]), .B1(\mem[208][3] ), .B2(n7459), 
        .Z(n1328) );
  OA22D0 U6749 ( .A1(n7460), .A2(prog_data[2]), .B1(\mem[208][2] ), .B2(n7459), 
        .Z(n1327) );
  OA22D0 U6750 ( .A1(n7460), .A2(prog_data[1]), .B1(\mem[208][1] ), .B2(n7459), 
        .Z(n1326) );
  OA22D0 U6751 ( .A1(n7460), .A2(prog_data[0]), .B1(\mem[208][0] ), .B2(n7459), 
        .Z(n1325) );
  NR2D0 U6752 ( .A1(n7531), .A2(n7489), .ZN(n7461) );
  INVD0 U6753 ( .I(n7461), .ZN(n7462) );
  OA22D0 U6754 ( .A1(n7462), .A2(prog_data[15]), .B1(\mem[209][15] ), .B2(
        n7461), .Z(n1324) );
  OA22D0 U6755 ( .A1(n7462), .A2(prog_data[14]), .B1(\mem[209][14] ), .B2(
        n7461), .Z(n1323) );
  OA22D0 U6756 ( .A1(n7462), .A2(prog_data[13]), .B1(\mem[209][13] ), .B2(
        n7461), .Z(n1322) );
  OA22D0 U6757 ( .A1(n7462), .A2(prog_data[12]), .B1(\mem[209][12] ), .B2(
        n7461), .Z(n1321) );
  OA22D0 U6758 ( .A1(n7462), .A2(prog_data[11]), .B1(\mem[209][11] ), .B2(
        n7461), .Z(n1320) );
  OA22D0 U6759 ( .A1(n7462), .A2(prog_data[10]), .B1(\mem[209][10] ), .B2(
        n7461), .Z(n1319) );
  OA22D0 U6760 ( .A1(n7462), .A2(prog_data[9]), .B1(\mem[209][9] ), .B2(n7461), 
        .Z(n1318) );
  OA22D0 U6761 ( .A1(n7462), .A2(prog_data[8]), .B1(\mem[209][8] ), .B2(n7461), 
        .Z(n1317) );
  OA22D0 U6762 ( .A1(n7462), .A2(prog_data[7]), .B1(\mem[209][7] ), .B2(n7461), 
        .Z(n1316) );
  OA22D0 U6763 ( .A1(n7462), .A2(prog_data[6]), .B1(\mem[209][6] ), .B2(n7461), 
        .Z(n1315) );
  OA22D0 U6764 ( .A1(n7462), .A2(prog_data[5]), .B1(\mem[209][5] ), .B2(n7461), 
        .Z(n1314) );
  OA22D0 U6765 ( .A1(n7462), .A2(prog_data[4]), .B1(\mem[209][4] ), .B2(n7461), 
        .Z(n1313) );
  OA22D0 U6766 ( .A1(n7462), .A2(prog_data[3]), .B1(\mem[209][3] ), .B2(n7461), 
        .Z(n1312) );
  OA22D0 U6767 ( .A1(n7462), .A2(prog_data[2]), .B1(\mem[209][2] ), .B2(n7461), 
        .Z(n1311) );
  OA22D0 U6768 ( .A1(n7462), .A2(prog_data[1]), .B1(\mem[209][1] ), .B2(n7461), 
        .Z(n1310) );
  OA22D0 U6769 ( .A1(n7462), .A2(prog_data[0]), .B1(\mem[209][0] ), .B2(n7461), 
        .Z(n1309) );
  NR2D0 U6770 ( .A1(n7534), .A2(n7489), .ZN(n7463) );
  INVD0 U6771 ( .I(n7463), .ZN(n7464) );
  OA22D0 U6772 ( .A1(n7464), .A2(prog_data[15]), .B1(\mem[210][15] ), .B2(
        n7463), .Z(n1308) );
  OA22D0 U6773 ( .A1(n7464), .A2(prog_data[14]), .B1(\mem[210][14] ), .B2(
        n7463), .Z(n1307) );
  OA22D0 U6774 ( .A1(n7464), .A2(prog_data[13]), .B1(\mem[210][13] ), .B2(
        n7463), .Z(n1306) );
  OA22D0 U6775 ( .A1(n7464), .A2(prog_data[12]), .B1(\mem[210][12] ), .B2(
        n7463), .Z(n1305) );
  OA22D0 U6776 ( .A1(n7464), .A2(prog_data[11]), .B1(\mem[210][11] ), .B2(
        n7463), .Z(n1304) );
  OA22D0 U6777 ( .A1(n7464), .A2(prog_data[10]), .B1(\mem[210][10] ), .B2(
        n7463), .Z(n1303) );
  OA22D0 U6778 ( .A1(n7464), .A2(prog_data[9]), .B1(\mem[210][9] ), .B2(n7463), 
        .Z(n1302) );
  OA22D0 U6779 ( .A1(n7464), .A2(prog_data[8]), .B1(\mem[210][8] ), .B2(n7463), 
        .Z(n1301) );
  OA22D0 U6780 ( .A1(n7464), .A2(prog_data[7]), .B1(\mem[210][7] ), .B2(n7463), 
        .Z(n1300) );
  OA22D0 U6781 ( .A1(n7464), .A2(prog_data[6]), .B1(\mem[210][6] ), .B2(n7463), 
        .Z(n1299) );
  OA22D0 U6782 ( .A1(n7464), .A2(prog_data[5]), .B1(\mem[210][5] ), .B2(n7463), 
        .Z(n1298) );
  OA22D0 U6783 ( .A1(n7464), .A2(prog_data[4]), .B1(\mem[210][4] ), .B2(n7463), 
        .Z(n1297) );
  OA22D0 U6784 ( .A1(n7464), .A2(prog_data[3]), .B1(\mem[210][3] ), .B2(n7463), 
        .Z(n1296) );
  OA22D0 U6785 ( .A1(n7464), .A2(prog_data[2]), .B1(\mem[210][2] ), .B2(n7463), 
        .Z(n1295) );
  OA22D0 U6786 ( .A1(n7464), .A2(prog_data[1]), .B1(\mem[210][1] ), .B2(n7463), 
        .Z(n1294) );
  OA22D0 U6787 ( .A1(n7464), .A2(prog_data[0]), .B1(\mem[210][0] ), .B2(n7463), 
        .Z(n1293) );
  INVD0 U6788 ( .I(n7465), .ZN(n7466) );
  OA22D0 U6789 ( .A1(n7466), .A2(prog_data[15]), .B1(\mem[211][15] ), .B2(
        n7465), .Z(n1292) );
  OA22D0 U6790 ( .A1(n7466), .A2(prog_data[14]), .B1(\mem[211][14] ), .B2(
        n7465), .Z(n1291) );
  OA22D0 U6791 ( .A1(n7466), .A2(prog_data[13]), .B1(\mem[211][13] ), .B2(
        n7465), .Z(n1290) );
  OA22D0 U6792 ( .A1(n7466), .A2(prog_data[12]), .B1(\mem[211][12] ), .B2(
        n7465), .Z(n1289) );
  OA22D0 U6793 ( .A1(n7466), .A2(prog_data[11]), .B1(\mem[211][11] ), .B2(
        n7465), .Z(n1288) );
  OA22D0 U6794 ( .A1(n7466), .A2(prog_data[10]), .B1(\mem[211][10] ), .B2(
        n7465), .Z(n1287) );
  OA22D0 U6795 ( .A1(n7466), .A2(prog_data[9]), .B1(\mem[211][9] ), .B2(n7465), 
        .Z(n1286) );
  OA22D0 U6796 ( .A1(n7466), .A2(prog_data[8]), .B1(\mem[211][8] ), .B2(n7465), 
        .Z(n1285) );
  OA22D0 U6797 ( .A1(n7466), .A2(prog_data[7]), .B1(\mem[211][7] ), .B2(n7465), 
        .Z(n1284) );
  OA22D0 U6798 ( .A1(n7466), .A2(prog_data[6]), .B1(\mem[211][6] ), .B2(n7465), 
        .Z(n1283) );
  OA22D0 U6799 ( .A1(n7466), .A2(prog_data[5]), .B1(\mem[211][5] ), .B2(n7465), 
        .Z(n1282) );
  OA22D0 U6800 ( .A1(n7466), .A2(prog_data[4]), .B1(\mem[211][4] ), .B2(n7465), 
        .Z(n1281) );
  OA22D0 U6801 ( .A1(n7466), .A2(prog_data[3]), .B1(\mem[211][3] ), .B2(n7465), 
        .Z(n1280) );
  OA22D0 U6802 ( .A1(n7466), .A2(prog_data[2]), .B1(\mem[211][2] ), .B2(n7465), 
        .Z(n1279) );
  OA22D0 U6803 ( .A1(n7466), .A2(prog_data[1]), .B1(\mem[211][1] ), .B2(n7465), 
        .Z(n1278) );
  OA22D0 U6804 ( .A1(n7466), .A2(prog_data[0]), .B1(\mem[211][0] ), .B2(n7465), 
        .Z(n1277) );
  NR2D0 U6805 ( .A1(n7540), .A2(n7489), .ZN(n7467) );
  INVD0 U6806 ( .I(n7467), .ZN(n7468) );
  OA22D0 U6807 ( .A1(n7468), .A2(prog_data[15]), .B1(\mem[212][15] ), .B2(
        n7467), .Z(n1276) );
  OA22D0 U6808 ( .A1(n7468), .A2(prog_data[14]), .B1(\mem[212][14] ), .B2(
        n7467), .Z(n1275) );
  OA22D0 U6809 ( .A1(n7468), .A2(prog_data[13]), .B1(\mem[212][13] ), .B2(
        n7467), .Z(n1274) );
  OA22D0 U6810 ( .A1(n7468), .A2(prog_data[12]), .B1(\mem[212][12] ), .B2(
        n7467), .Z(n1273) );
  OA22D0 U6811 ( .A1(n7468), .A2(prog_data[11]), .B1(\mem[212][11] ), .B2(
        n7467), .Z(n1272) );
  OA22D0 U6812 ( .A1(n7468), .A2(prog_data[10]), .B1(\mem[212][10] ), .B2(
        n7467), .Z(n1271) );
  OA22D0 U6813 ( .A1(n7468), .A2(prog_data[9]), .B1(\mem[212][9] ), .B2(n7467), 
        .Z(n1270) );
  OA22D0 U6814 ( .A1(n7468), .A2(prog_data[8]), .B1(\mem[212][8] ), .B2(n7467), 
        .Z(n1269) );
  OA22D0 U6815 ( .A1(n7468), .A2(prog_data[7]), .B1(\mem[212][7] ), .B2(n7467), 
        .Z(n1268) );
  OA22D0 U6816 ( .A1(n7468), .A2(prog_data[6]), .B1(\mem[212][6] ), .B2(n7467), 
        .Z(n1267) );
  OA22D0 U6817 ( .A1(n7468), .A2(prog_data[5]), .B1(\mem[212][5] ), .B2(n7467), 
        .Z(n1266) );
  OA22D0 U6818 ( .A1(n7468), .A2(prog_data[4]), .B1(\mem[212][4] ), .B2(n7467), 
        .Z(n1265) );
  OA22D0 U6819 ( .A1(n7468), .A2(prog_data[3]), .B1(\mem[212][3] ), .B2(n7467), 
        .Z(n1264) );
  OA22D0 U6820 ( .A1(n7468), .A2(prog_data[2]), .B1(\mem[212][2] ), .B2(n7467), 
        .Z(n1263) );
  OA22D0 U6821 ( .A1(n7468), .A2(prog_data[1]), .B1(\mem[212][1] ), .B2(n7467), 
        .Z(n1262) );
  OA22D0 U6822 ( .A1(n7468), .A2(prog_data[0]), .B1(\mem[212][0] ), .B2(n7467), 
        .Z(n1261) );
  NR2D0 U6823 ( .A1(n7543), .A2(n7489), .ZN(n7469) );
  INVD0 U6824 ( .I(n7469), .ZN(n7470) );
  OA22D0 U6825 ( .A1(n7470), .A2(prog_data[15]), .B1(\mem[213][15] ), .B2(
        n7469), .Z(n1260) );
  OA22D0 U6826 ( .A1(n7470), .A2(prog_data[14]), .B1(\mem[213][14] ), .B2(
        n7469), .Z(n1259) );
  OA22D0 U6827 ( .A1(n7470), .A2(prog_data[13]), .B1(\mem[213][13] ), .B2(
        n7469), .Z(n1258) );
  OA22D0 U6828 ( .A1(n7470), .A2(prog_data[12]), .B1(\mem[213][12] ), .B2(
        n7469), .Z(n1257) );
  OA22D0 U6829 ( .A1(n7470), .A2(prog_data[11]), .B1(\mem[213][11] ), .B2(
        n7469), .Z(n1256) );
  OA22D0 U6830 ( .A1(n7470), .A2(prog_data[10]), .B1(\mem[213][10] ), .B2(
        n7469), .Z(n1255) );
  OA22D0 U6831 ( .A1(n7470), .A2(prog_data[9]), .B1(\mem[213][9] ), .B2(n7469), 
        .Z(n1254) );
  OA22D0 U6832 ( .A1(n7470), .A2(prog_data[8]), .B1(\mem[213][8] ), .B2(n7469), 
        .Z(n1253) );
  OA22D0 U6833 ( .A1(n7470), .A2(prog_data[7]), .B1(\mem[213][7] ), .B2(n7469), 
        .Z(n1252) );
  OA22D0 U6834 ( .A1(n7470), .A2(prog_data[6]), .B1(\mem[213][6] ), .B2(n7469), 
        .Z(n1251) );
  OA22D0 U6835 ( .A1(n7470), .A2(prog_data[5]), .B1(\mem[213][5] ), .B2(n7469), 
        .Z(n1250) );
  OA22D0 U6836 ( .A1(n7470), .A2(prog_data[4]), .B1(\mem[213][4] ), .B2(n7469), 
        .Z(n1249) );
  OA22D0 U6837 ( .A1(n7470), .A2(prog_data[3]), .B1(\mem[213][3] ), .B2(n7469), 
        .Z(n1248) );
  OA22D0 U6838 ( .A1(n7470), .A2(prog_data[2]), .B1(\mem[213][2] ), .B2(n7469), 
        .Z(n1247) );
  OA22D0 U6839 ( .A1(n7470), .A2(prog_data[1]), .B1(\mem[213][1] ), .B2(n7469), 
        .Z(n1246) );
  OA22D0 U6840 ( .A1(n7470), .A2(prog_data[0]), .B1(\mem[213][0] ), .B2(n7469), 
        .Z(n1245) );
  NR2D0 U6841 ( .A1(n7546), .A2(n7489), .ZN(n7471) );
  INVD0 U6842 ( .I(n7471), .ZN(n7472) );
  OA22D0 U6843 ( .A1(n7472), .A2(prog_data[15]), .B1(\mem[214][15] ), .B2(
        n7471), .Z(n1244) );
  OA22D0 U6844 ( .A1(n7472), .A2(prog_data[14]), .B1(\mem[214][14] ), .B2(
        n7471), .Z(n1243) );
  OA22D0 U6845 ( .A1(n7472), .A2(prog_data[13]), .B1(\mem[214][13] ), .B2(
        n7471), .Z(n1242) );
  OA22D0 U6846 ( .A1(n7472), .A2(prog_data[12]), .B1(\mem[214][12] ), .B2(
        n7471), .Z(n1241) );
  OA22D0 U6847 ( .A1(n7472), .A2(prog_data[11]), .B1(\mem[214][11] ), .B2(
        n7471), .Z(n1240) );
  OA22D0 U6848 ( .A1(n7472), .A2(prog_data[10]), .B1(\mem[214][10] ), .B2(
        n7471), .Z(n1239) );
  OA22D0 U6849 ( .A1(n7472), .A2(prog_data[9]), .B1(\mem[214][9] ), .B2(n7471), 
        .Z(n1238) );
  OA22D0 U6850 ( .A1(n7472), .A2(prog_data[8]), .B1(\mem[214][8] ), .B2(n7471), 
        .Z(n1237) );
  OA22D0 U6851 ( .A1(n7472), .A2(prog_data[7]), .B1(\mem[214][7] ), .B2(n7471), 
        .Z(n1236) );
  OA22D0 U6852 ( .A1(n7472), .A2(prog_data[6]), .B1(\mem[214][6] ), .B2(n7471), 
        .Z(n1235) );
  OA22D0 U6853 ( .A1(n7472), .A2(prog_data[5]), .B1(\mem[214][5] ), .B2(n7471), 
        .Z(n1234) );
  OA22D0 U6854 ( .A1(n7472), .A2(prog_data[4]), .B1(\mem[214][4] ), .B2(n7471), 
        .Z(n1233) );
  OA22D0 U6855 ( .A1(n7472), .A2(prog_data[3]), .B1(\mem[214][3] ), .B2(n7471), 
        .Z(n1232) );
  OA22D0 U6856 ( .A1(n7472), .A2(prog_data[2]), .B1(\mem[214][2] ), .B2(n7471), 
        .Z(n1231) );
  OA22D0 U6857 ( .A1(n7472), .A2(prog_data[1]), .B1(\mem[214][1] ), .B2(n7471), 
        .Z(n1230) );
  OA22D0 U6858 ( .A1(n7472), .A2(prog_data[0]), .B1(\mem[214][0] ), .B2(n7471), 
        .Z(n1229) );
  NR2D0 U6859 ( .A1(n7549), .A2(n7489), .ZN(n7473) );
  INVD0 U6860 ( .I(n7473), .ZN(n7474) );
  OA22D0 U6861 ( .A1(n7474), .A2(prog_data[15]), .B1(\mem[215][15] ), .B2(
        n7473), .Z(n1228) );
  OA22D0 U6862 ( .A1(n7474), .A2(prog_data[14]), .B1(\mem[215][14] ), .B2(
        n7473), .Z(n1227) );
  OA22D0 U6863 ( .A1(n7474), .A2(prog_data[13]), .B1(\mem[215][13] ), .B2(
        n7473), .Z(n1226) );
  OA22D0 U6864 ( .A1(n7474), .A2(prog_data[12]), .B1(\mem[215][12] ), .B2(
        n7473), .Z(n1225) );
  OA22D0 U6865 ( .A1(n7474), .A2(prog_data[11]), .B1(\mem[215][11] ), .B2(
        n7473), .Z(n1224) );
  OA22D0 U6866 ( .A1(n7474), .A2(prog_data[10]), .B1(\mem[215][10] ), .B2(
        n7473), .Z(n1223) );
  OA22D0 U6867 ( .A1(n7474), .A2(prog_data[9]), .B1(\mem[215][9] ), .B2(n7473), 
        .Z(n1222) );
  OA22D0 U6868 ( .A1(n7474), .A2(prog_data[8]), .B1(\mem[215][8] ), .B2(n7473), 
        .Z(n1221) );
  OA22D0 U6869 ( .A1(n7474), .A2(prog_data[7]), .B1(\mem[215][7] ), .B2(n7473), 
        .Z(n1220) );
  OA22D0 U6870 ( .A1(n7474), .A2(prog_data[6]), .B1(\mem[215][6] ), .B2(n7473), 
        .Z(n1219) );
  OA22D0 U6871 ( .A1(n7474), .A2(prog_data[5]), .B1(\mem[215][5] ), .B2(n7473), 
        .Z(n1218) );
  OA22D0 U6872 ( .A1(n7474), .A2(prog_data[4]), .B1(\mem[215][4] ), .B2(n7473), 
        .Z(n1217) );
  OA22D0 U6873 ( .A1(n7474), .A2(prog_data[3]), .B1(\mem[215][3] ), .B2(n7473), 
        .Z(n1216) );
  OA22D0 U6874 ( .A1(n7474), .A2(prog_data[2]), .B1(\mem[215][2] ), .B2(n7473), 
        .Z(n1215) );
  OA22D0 U6875 ( .A1(n7474), .A2(prog_data[1]), .B1(\mem[215][1] ), .B2(n7473), 
        .Z(n1214) );
  OA22D0 U6876 ( .A1(n7474), .A2(prog_data[0]), .B1(\mem[215][0] ), .B2(n7473), 
        .Z(n1213) );
  NR2D0 U6877 ( .A1(n7552), .A2(n7489), .ZN(n7475) );
  INVD0 U6878 ( .I(n7475), .ZN(n7476) );
  OA22D0 U6879 ( .A1(n7476), .A2(prog_data[15]), .B1(\mem[216][15] ), .B2(
        n7475), .Z(n1212) );
  OA22D0 U6880 ( .A1(n7476), .A2(prog_data[14]), .B1(\mem[216][14] ), .B2(
        n7475), .Z(n1211) );
  OA22D0 U6881 ( .A1(n7476), .A2(prog_data[13]), .B1(\mem[216][13] ), .B2(
        n7475), .Z(n1210) );
  OA22D0 U6882 ( .A1(n7476), .A2(prog_data[12]), .B1(\mem[216][12] ), .B2(
        n7475), .Z(n1209) );
  OA22D0 U6883 ( .A1(n7476), .A2(prog_data[11]), .B1(\mem[216][11] ), .B2(
        n7475), .Z(n1208) );
  OA22D0 U6884 ( .A1(n7476), .A2(prog_data[10]), .B1(\mem[216][10] ), .B2(
        n7475), .Z(n1207) );
  OA22D0 U6885 ( .A1(n7476), .A2(prog_data[9]), .B1(\mem[216][9] ), .B2(n7475), 
        .Z(n1206) );
  OA22D0 U6886 ( .A1(n7476), .A2(prog_data[8]), .B1(\mem[216][8] ), .B2(n7475), 
        .Z(n1205) );
  OA22D0 U6887 ( .A1(n7476), .A2(prog_data[7]), .B1(\mem[216][7] ), .B2(n7475), 
        .Z(n1204) );
  OA22D0 U6888 ( .A1(n7476), .A2(prog_data[6]), .B1(\mem[216][6] ), .B2(n7475), 
        .Z(n1203) );
  OA22D0 U6889 ( .A1(n7476), .A2(prog_data[5]), .B1(\mem[216][5] ), .B2(n7475), 
        .Z(n1202) );
  OA22D0 U6890 ( .A1(n7476), .A2(prog_data[4]), .B1(\mem[216][4] ), .B2(n7475), 
        .Z(n1201) );
  OA22D0 U6891 ( .A1(n7476), .A2(prog_data[3]), .B1(\mem[216][3] ), .B2(n7475), 
        .Z(n1200) );
  OA22D0 U6892 ( .A1(n7476), .A2(prog_data[2]), .B1(\mem[216][2] ), .B2(n7475), 
        .Z(n1199) );
  OA22D0 U6893 ( .A1(n7476), .A2(prog_data[1]), .B1(\mem[216][1] ), .B2(n7475), 
        .Z(n1198) );
  OA22D0 U6894 ( .A1(n7476), .A2(prog_data[0]), .B1(\mem[216][0] ), .B2(n7475), 
        .Z(n1197) );
  NR2D0 U6895 ( .A1(n7555), .A2(n7489), .ZN(n7477) );
  INVD0 U6896 ( .I(n7477), .ZN(n7478) );
  OA22D0 U6897 ( .A1(n7478), .A2(prog_data[15]), .B1(\mem[217][15] ), .B2(
        n7477), .Z(n1196) );
  OA22D0 U6898 ( .A1(n7478), .A2(prog_data[14]), .B1(\mem[217][14] ), .B2(
        n7477), .Z(n1195) );
  OA22D0 U6899 ( .A1(n7478), .A2(prog_data[13]), .B1(\mem[217][13] ), .B2(
        n7477), .Z(n1194) );
  OA22D0 U6900 ( .A1(n7478), .A2(prog_data[12]), .B1(\mem[217][12] ), .B2(
        n7477), .Z(n1193) );
  OA22D0 U6901 ( .A1(n7478), .A2(prog_data[11]), .B1(\mem[217][11] ), .B2(
        n7477), .Z(n1192) );
  OA22D0 U6902 ( .A1(n7478), .A2(prog_data[10]), .B1(\mem[217][10] ), .B2(
        n7477), .Z(n1191) );
  OA22D0 U6903 ( .A1(n7478), .A2(prog_data[9]), .B1(\mem[217][9] ), .B2(n7477), 
        .Z(n1190) );
  OA22D0 U6904 ( .A1(n7478), .A2(prog_data[8]), .B1(\mem[217][8] ), .B2(n7477), 
        .Z(n1189) );
  OA22D0 U6905 ( .A1(n7478), .A2(prog_data[7]), .B1(\mem[217][7] ), .B2(n7477), 
        .Z(n1188) );
  OA22D0 U6906 ( .A1(n7478), .A2(prog_data[6]), .B1(\mem[217][6] ), .B2(n7477), 
        .Z(n1187) );
  OA22D0 U6907 ( .A1(n7478), .A2(prog_data[5]), .B1(\mem[217][5] ), .B2(n7477), 
        .Z(n1186) );
  OA22D0 U6908 ( .A1(n7478), .A2(prog_data[4]), .B1(\mem[217][4] ), .B2(n7477), 
        .Z(n1185) );
  OA22D0 U6909 ( .A1(n7478), .A2(prog_data[3]), .B1(\mem[217][3] ), .B2(n7477), 
        .Z(n1184) );
  OA22D0 U6910 ( .A1(n7478), .A2(prog_data[2]), .B1(\mem[217][2] ), .B2(n7477), 
        .Z(n1183) );
  OA22D0 U6911 ( .A1(n7478), .A2(prog_data[1]), .B1(\mem[217][1] ), .B2(n7477), 
        .Z(n1182) );
  OA22D0 U6912 ( .A1(n7478), .A2(prog_data[0]), .B1(\mem[217][0] ), .B2(n7477), 
        .Z(n1181) );
  NR2D0 U6913 ( .A1(n7558), .A2(n7489), .ZN(n7479) );
  INVD0 U6914 ( .I(n7479), .ZN(n7480) );
  OA22D0 U6915 ( .A1(n7480), .A2(prog_data[15]), .B1(\mem[218][15] ), .B2(
        n7479), .Z(n1180) );
  OA22D0 U6916 ( .A1(n7480), .A2(prog_data[14]), .B1(\mem[218][14] ), .B2(
        n7479), .Z(n1179) );
  OA22D0 U6917 ( .A1(n7480), .A2(prog_data[13]), .B1(\mem[218][13] ), .B2(
        n7479), .Z(n1178) );
  OA22D0 U6918 ( .A1(n7480), .A2(prog_data[12]), .B1(\mem[218][12] ), .B2(
        n7479), .Z(n1177) );
  OA22D0 U6919 ( .A1(n7480), .A2(prog_data[11]), .B1(\mem[218][11] ), .B2(
        n7479), .Z(n1176) );
  OA22D0 U6920 ( .A1(n7480), .A2(prog_data[10]), .B1(\mem[218][10] ), .B2(
        n7479), .Z(n1175) );
  OA22D0 U6921 ( .A1(n7480), .A2(prog_data[9]), .B1(\mem[218][9] ), .B2(n7479), 
        .Z(n1174) );
  OA22D0 U6922 ( .A1(n7480), .A2(prog_data[8]), .B1(\mem[218][8] ), .B2(n7479), 
        .Z(n1173) );
  OA22D0 U6923 ( .A1(n7480), .A2(prog_data[7]), .B1(\mem[218][7] ), .B2(n7479), 
        .Z(n1172) );
  OA22D0 U6924 ( .A1(n7480), .A2(prog_data[6]), .B1(\mem[218][6] ), .B2(n7479), 
        .Z(n1171) );
  OA22D0 U6925 ( .A1(n7480), .A2(prog_data[5]), .B1(\mem[218][5] ), .B2(n7479), 
        .Z(n1170) );
  OA22D0 U6926 ( .A1(n7480), .A2(prog_data[4]), .B1(\mem[218][4] ), .B2(n7479), 
        .Z(n1169) );
  OA22D0 U6927 ( .A1(n7480), .A2(prog_data[3]), .B1(\mem[218][3] ), .B2(n7479), 
        .Z(n1168) );
  OA22D0 U6928 ( .A1(n7480), .A2(prog_data[2]), .B1(\mem[218][2] ), .B2(n7479), 
        .Z(n1167) );
  OA22D0 U6929 ( .A1(n7480), .A2(prog_data[1]), .B1(\mem[218][1] ), .B2(n7479), 
        .Z(n1166) );
  OA22D0 U6930 ( .A1(n7480), .A2(prog_data[0]), .B1(\mem[218][0] ), .B2(n7479), 
        .Z(n1165) );
  NR2D0 U6931 ( .A1(n7561), .A2(n7489), .ZN(n7481) );
  OA22D0 U6932 ( .A1(n7482), .A2(prog_data[15]), .B1(\mem[219][15] ), .B2(
        n7481), .Z(n1164) );
  OA22D0 U6933 ( .A1(n7482), .A2(prog_data[14]), .B1(\mem[219][14] ), .B2(
        n7481), .Z(n1163) );
  OA22D0 U6934 ( .A1(n7482), .A2(prog_data[13]), .B1(\mem[219][13] ), .B2(
        n7481), .Z(n1162) );
  OA22D0 U6935 ( .A1(n7482), .A2(prog_data[12]), .B1(\mem[219][12] ), .B2(
        n7481), .Z(n1161) );
  OA22D0 U6936 ( .A1(n7482), .A2(prog_data[11]), .B1(\mem[219][11] ), .B2(
        n7481), .Z(n1160) );
  OA22D0 U6937 ( .A1(n7482), .A2(prog_data[10]), .B1(\mem[219][10] ), .B2(
        n7481), .Z(n1159) );
  OA22D0 U6938 ( .A1(n7482), .A2(prog_data[9]), .B1(\mem[219][9] ), .B2(n7481), 
        .Z(n1158) );
  OA22D0 U6939 ( .A1(n7482), .A2(prog_data[8]), .B1(\mem[219][8] ), .B2(n7481), 
        .Z(n1157) );
  OA22D0 U6940 ( .A1(n7482), .A2(prog_data[7]), .B1(\mem[219][7] ), .B2(n7481), 
        .Z(n1156) );
  OA22D0 U6941 ( .A1(n7482), .A2(prog_data[6]), .B1(\mem[219][6] ), .B2(n7481), 
        .Z(n1155) );
  OA22D0 U6942 ( .A1(n7482), .A2(prog_data[5]), .B1(\mem[219][5] ), .B2(n7481), 
        .Z(n1154) );
  OA22D0 U6943 ( .A1(n7482), .A2(prog_data[4]), .B1(\mem[219][4] ), .B2(n7481), 
        .Z(n1153) );
  OA22D0 U6944 ( .A1(n7482), .A2(prog_data[3]), .B1(\mem[219][3] ), .B2(n7481), 
        .Z(n1152) );
  OA22D0 U6945 ( .A1(n7482), .A2(prog_data[2]), .B1(\mem[219][2] ), .B2(n7481), 
        .Z(n1151) );
  OA22D0 U6946 ( .A1(n7482), .A2(prog_data[1]), .B1(\mem[219][1] ), .B2(n7481), 
        .Z(n1150) );
  OA22D0 U6947 ( .A1(n7482), .A2(prog_data[0]), .B1(\mem[219][0] ), .B2(n7481), 
        .Z(n1149) );
  NR2D0 U6948 ( .A1(n7564), .A2(n7489), .ZN(n7483) );
  INVD0 U6949 ( .I(n7483), .ZN(n7484) );
  OA22D0 U6950 ( .A1(n7484), .A2(prog_data[15]), .B1(\mem[220][15] ), .B2(
        n7483), .Z(n1148) );
  OA22D0 U6951 ( .A1(n7484), .A2(prog_data[14]), .B1(\mem[220][14] ), .B2(
        n7483), .Z(n1147) );
  OA22D0 U6952 ( .A1(n7484), .A2(prog_data[13]), .B1(\mem[220][13] ), .B2(
        n7483), .Z(n1146) );
  OA22D0 U6953 ( .A1(n7484), .A2(prog_data[12]), .B1(\mem[220][12] ), .B2(
        n7483), .Z(n1145) );
  OA22D0 U6954 ( .A1(n7484), .A2(prog_data[11]), .B1(\mem[220][11] ), .B2(
        n7483), .Z(n1144) );
  OA22D0 U6955 ( .A1(n7484), .A2(prog_data[10]), .B1(\mem[220][10] ), .B2(
        n7483), .Z(n1143) );
  OA22D0 U6956 ( .A1(n7484), .A2(prog_data[9]), .B1(\mem[220][9] ), .B2(n7483), 
        .Z(n1142) );
  OA22D0 U6957 ( .A1(n7484), .A2(prog_data[8]), .B1(\mem[220][8] ), .B2(n7483), 
        .Z(n1141) );
  OA22D0 U6958 ( .A1(n7484), .A2(prog_data[7]), .B1(\mem[220][7] ), .B2(n7483), 
        .Z(n1140) );
  OA22D0 U6959 ( .A1(n7484), .A2(prog_data[6]), .B1(\mem[220][6] ), .B2(n7483), 
        .Z(n1139) );
  OA22D0 U6960 ( .A1(n7484), .A2(prog_data[5]), .B1(\mem[220][5] ), .B2(n7483), 
        .Z(n1138) );
  OA22D0 U6961 ( .A1(n7484), .A2(prog_data[4]), .B1(\mem[220][4] ), .B2(n7483), 
        .Z(n1137) );
  OA22D0 U6962 ( .A1(n7484), .A2(prog_data[3]), .B1(\mem[220][3] ), .B2(n7483), 
        .Z(n1136) );
  OA22D0 U6963 ( .A1(n7484), .A2(prog_data[2]), .B1(\mem[220][2] ), .B2(n7483), 
        .Z(n1135) );
  OA22D0 U6964 ( .A1(n7484), .A2(prog_data[1]), .B1(\mem[220][1] ), .B2(n7483), 
        .Z(n1134) );
  OA22D0 U6965 ( .A1(n7484), .A2(prog_data[0]), .B1(\mem[220][0] ), .B2(n7483), 
        .Z(n1133) );
  NR2D0 U6966 ( .A1(n7567), .A2(n7489), .ZN(n7485) );
  INVD0 U6967 ( .I(n7485), .ZN(n7486) );
  OA22D0 U6968 ( .A1(n7486), .A2(prog_data[15]), .B1(\mem[221][15] ), .B2(
        n7485), .Z(n1132) );
  OA22D0 U6969 ( .A1(n7486), .A2(prog_data[14]), .B1(\mem[221][14] ), .B2(
        n7485), .Z(n1131) );
  OA22D0 U6970 ( .A1(n7486), .A2(prog_data[13]), .B1(\mem[221][13] ), .B2(
        n7485), .Z(n1130) );
  OA22D0 U6971 ( .A1(n7486), .A2(prog_data[12]), .B1(\mem[221][12] ), .B2(
        n7485), .Z(n1129) );
  OA22D0 U6972 ( .A1(n7486), .A2(prog_data[11]), .B1(\mem[221][11] ), .B2(
        n7485), .Z(n1128) );
  OA22D0 U6973 ( .A1(n7486), .A2(prog_data[10]), .B1(\mem[221][10] ), .B2(
        n7485), .Z(n1127) );
  OA22D0 U6974 ( .A1(n7486), .A2(prog_data[9]), .B1(\mem[221][9] ), .B2(n7485), 
        .Z(n1126) );
  OA22D0 U6975 ( .A1(n7486), .A2(prog_data[8]), .B1(\mem[221][8] ), .B2(n7485), 
        .Z(n1125) );
  OA22D0 U6976 ( .A1(n7486), .A2(prog_data[7]), .B1(\mem[221][7] ), .B2(n7485), 
        .Z(n1124) );
  OA22D0 U6977 ( .A1(n7486), .A2(prog_data[6]), .B1(\mem[221][6] ), .B2(n7485), 
        .Z(n1123) );
  OA22D0 U6978 ( .A1(n7486), .A2(prog_data[5]), .B1(\mem[221][5] ), .B2(n7485), 
        .Z(n1122) );
  OA22D0 U6979 ( .A1(n7486), .A2(prog_data[4]), .B1(\mem[221][4] ), .B2(n7485), 
        .Z(n1121) );
  OA22D0 U6980 ( .A1(n7486), .A2(prog_data[3]), .B1(\mem[221][3] ), .B2(n7485), 
        .Z(n1120) );
  OA22D0 U6981 ( .A1(n7486), .A2(prog_data[2]), .B1(\mem[221][2] ), .B2(n7485), 
        .Z(n1119) );
  OA22D0 U6982 ( .A1(n7486), .A2(prog_data[1]), .B1(\mem[221][1] ), .B2(n7485), 
        .Z(n1118) );
  OA22D0 U6983 ( .A1(n7486), .A2(prog_data[0]), .B1(\mem[221][0] ), .B2(n7485), 
        .Z(n1117) );
  NR2D0 U6984 ( .A1(n7570), .A2(n7489), .ZN(n7487) );
  INVD0 U6985 ( .I(n7487), .ZN(n7488) );
  OA22D0 U6986 ( .A1(n7488), .A2(prog_data[15]), .B1(\mem[222][15] ), .B2(
        n7487), .Z(n1116) );
  OA22D0 U6987 ( .A1(n7488), .A2(prog_data[14]), .B1(\mem[222][14] ), .B2(
        n7487), .Z(n1115) );
  OA22D0 U6988 ( .A1(n7488), .A2(prog_data[13]), .B1(\mem[222][13] ), .B2(
        n7487), .Z(n1114) );
  OA22D0 U6989 ( .A1(n7488), .A2(prog_data[12]), .B1(\mem[222][12] ), .B2(
        n7487), .Z(n1113) );
  OA22D0 U6990 ( .A1(n7488), .A2(prog_data[11]), .B1(\mem[222][11] ), .B2(
        n7487), .Z(n1112) );
  OA22D0 U6991 ( .A1(n7488), .A2(prog_data[10]), .B1(\mem[222][10] ), .B2(
        n7487), .Z(n1111) );
  OA22D0 U6992 ( .A1(n7488), .A2(prog_data[9]), .B1(\mem[222][9] ), .B2(n7487), 
        .Z(n1110) );
  OA22D0 U6993 ( .A1(n7488), .A2(prog_data[8]), .B1(\mem[222][8] ), .B2(n7487), 
        .Z(n1109) );
  OA22D0 U6994 ( .A1(n7488), .A2(prog_data[7]), .B1(\mem[222][7] ), .B2(n7487), 
        .Z(n1108) );
  OA22D0 U6995 ( .A1(n7488), .A2(prog_data[6]), .B1(\mem[222][6] ), .B2(n7487), 
        .Z(n1107) );
  OA22D0 U6996 ( .A1(n7488), .A2(prog_data[5]), .B1(\mem[222][5] ), .B2(n7487), 
        .Z(n1106) );
  OA22D0 U6997 ( .A1(n7488), .A2(prog_data[4]), .B1(\mem[222][4] ), .B2(n7487), 
        .Z(n1105) );
  OA22D0 U6998 ( .A1(n7488), .A2(prog_data[3]), .B1(\mem[222][3] ), .B2(n7487), 
        .Z(n1104) );
  OA22D0 U6999 ( .A1(n7488), .A2(prog_data[2]), .B1(\mem[222][2] ), .B2(n7487), 
        .Z(n1103) );
  OA22D0 U7000 ( .A1(n7488), .A2(prog_data[1]), .B1(\mem[222][1] ), .B2(n7487), 
        .Z(n1102) );
  OA22D0 U7001 ( .A1(n7488), .A2(prog_data[0]), .B1(\mem[222][0] ), .B2(n7487), 
        .Z(n1101) );
  NR2D0 U7002 ( .A1(n7574), .A2(n7489), .ZN(n7490) );
  INVD0 U7003 ( .I(n7490), .ZN(n7491) );
  OA22D0 U7004 ( .A1(n7491), .A2(prog_data[15]), .B1(\mem[223][15] ), .B2(
        n7490), .Z(n1100) );
  OA22D0 U7005 ( .A1(n7491), .A2(prog_data[14]), .B1(\mem[223][14] ), .B2(
        n7490), .Z(n1099) );
  OA22D0 U7006 ( .A1(n7491), .A2(prog_data[13]), .B1(\mem[223][13] ), .B2(
        n7490), .Z(n1098) );
  OA22D0 U7007 ( .A1(n7491), .A2(prog_data[12]), .B1(\mem[223][12] ), .B2(
        n7490), .Z(n1097) );
  OA22D0 U7008 ( .A1(n7491), .A2(prog_data[11]), .B1(\mem[223][11] ), .B2(
        n7490), .Z(n1096) );
  OA22D0 U7009 ( .A1(n7491), .A2(prog_data[10]), .B1(\mem[223][10] ), .B2(
        n7490), .Z(n1095) );
  OA22D0 U7010 ( .A1(n7491), .A2(prog_data[9]), .B1(\mem[223][9] ), .B2(n7490), 
        .Z(n1094) );
  OA22D0 U7011 ( .A1(n7491), .A2(prog_data[8]), .B1(\mem[223][8] ), .B2(n7490), 
        .Z(n1093) );
  OA22D0 U7012 ( .A1(n7491), .A2(prog_data[7]), .B1(\mem[223][7] ), .B2(n7490), 
        .Z(n1092) );
  OA22D0 U7013 ( .A1(n7491), .A2(prog_data[6]), .B1(\mem[223][6] ), .B2(n7490), 
        .Z(n1091) );
  OA22D0 U7014 ( .A1(n7491), .A2(prog_data[5]), .B1(\mem[223][5] ), .B2(n7490), 
        .Z(n1090) );
  OA22D0 U7015 ( .A1(n7491), .A2(prog_data[4]), .B1(\mem[223][4] ), .B2(n7490), 
        .Z(n1089) );
  OA22D0 U7016 ( .A1(n7491), .A2(prog_data[3]), .B1(\mem[223][3] ), .B2(n7490), 
        .Z(n1088) );
  OA22D0 U7017 ( .A1(n7491), .A2(prog_data[2]), .B1(\mem[223][2] ), .B2(n7490), 
        .Z(n1087) );
  OA22D0 U7018 ( .A1(n7491), .A2(prog_data[1]), .B1(\mem[223][1] ), .B2(n7490), 
        .Z(n1086) );
  OA22D0 U7019 ( .A1(n7491), .A2(prog_data[0]), .B1(\mem[223][0] ), .B2(n7490), 
        .Z(n1085) );
  IND3D0 U7020 ( .A1(n7527), .B1(prog_addr[6]), .B2(n7492), .ZN(n7523) );
  NR2D0 U7021 ( .A1(n7528), .A2(n7523), .ZN(n7493) );
  INVD0 U7022 ( .I(n7493), .ZN(n7494) );
  OA22D0 U7023 ( .A1(n7494), .A2(prog_data[15]), .B1(\mem[224][15] ), .B2(
        n7493), .Z(n1084) );
  OA22D0 U7024 ( .A1(n7494), .A2(prog_data[14]), .B1(\mem[224][14] ), .B2(
        n7493), .Z(n1083) );
  OA22D0 U7025 ( .A1(n7494), .A2(prog_data[13]), .B1(\mem[224][13] ), .B2(
        n7493), .Z(n1082) );
  OA22D0 U7026 ( .A1(n7494), .A2(prog_data[12]), .B1(\mem[224][12] ), .B2(
        n7493), .Z(n1081) );
  OA22D0 U7027 ( .A1(n7494), .A2(prog_data[11]), .B1(\mem[224][11] ), .B2(
        n7493), .Z(n1080) );
  OA22D0 U7028 ( .A1(n7494), .A2(prog_data[10]), .B1(\mem[224][10] ), .B2(
        n7493), .Z(n1079) );
  OA22D0 U7029 ( .A1(n7494), .A2(prog_data[9]), .B1(\mem[224][9] ), .B2(n7493), 
        .Z(n1078) );
  OA22D0 U7030 ( .A1(n7494), .A2(prog_data[8]), .B1(\mem[224][8] ), .B2(n7493), 
        .Z(n1077) );
  OA22D0 U7031 ( .A1(n7494), .A2(prog_data[7]), .B1(\mem[224][7] ), .B2(n7493), 
        .Z(n1076) );
  OA22D0 U7032 ( .A1(n7494), .A2(prog_data[6]), .B1(\mem[224][6] ), .B2(n7493), 
        .Z(n1075) );
  OA22D0 U7033 ( .A1(n7494), .A2(prog_data[5]), .B1(\mem[224][5] ), .B2(n7493), 
        .Z(n1074) );
  OA22D0 U7034 ( .A1(n7494), .A2(prog_data[4]), .B1(\mem[224][4] ), .B2(n7493), 
        .Z(n1073) );
  OA22D0 U7035 ( .A1(n7494), .A2(prog_data[3]), .B1(\mem[224][3] ), .B2(n7493), 
        .Z(n1072) );
  OA22D0 U7036 ( .A1(n7494), .A2(prog_data[2]), .B1(\mem[224][2] ), .B2(n7493), 
        .Z(n1071) );
  OA22D0 U7037 ( .A1(n7494), .A2(prog_data[1]), .B1(\mem[224][1] ), .B2(n7493), 
        .Z(n1070) );
  OA22D0 U7038 ( .A1(n7494), .A2(prog_data[0]), .B1(\mem[224][0] ), .B2(n7493), 
        .Z(n1069) );
  NR2D0 U7039 ( .A1(n7531), .A2(n7523), .ZN(n7495) );
  INVD0 U7040 ( .I(n7495), .ZN(n7496) );
  OA22D0 U7041 ( .A1(n7496), .A2(prog_data[15]), .B1(\mem[225][15] ), .B2(
        n7495), .Z(n1068) );
  OA22D0 U7042 ( .A1(n7496), .A2(prog_data[14]), .B1(\mem[225][14] ), .B2(
        n7495), .Z(n1067) );
  OA22D0 U7043 ( .A1(n7496), .A2(prog_data[13]), .B1(\mem[225][13] ), .B2(
        n7495), .Z(n1066) );
  OA22D0 U7044 ( .A1(n7496), .A2(prog_data[12]), .B1(\mem[225][12] ), .B2(
        n7495), .Z(n1065) );
  OA22D0 U7045 ( .A1(n7496), .A2(prog_data[11]), .B1(\mem[225][11] ), .B2(
        n7495), .Z(n1064) );
  OA22D0 U7046 ( .A1(n7496), .A2(prog_data[10]), .B1(\mem[225][10] ), .B2(
        n7495), .Z(n1063) );
  OA22D0 U7047 ( .A1(n7496), .A2(prog_data[9]), .B1(\mem[225][9] ), .B2(n7495), 
        .Z(n1062) );
  OA22D0 U7048 ( .A1(n7496), .A2(prog_data[8]), .B1(\mem[225][8] ), .B2(n7495), 
        .Z(n1061) );
  OA22D0 U7049 ( .A1(n7496), .A2(prog_data[7]), .B1(\mem[225][7] ), .B2(n7495), 
        .Z(n1060) );
  OA22D0 U7050 ( .A1(n7496), .A2(prog_data[6]), .B1(\mem[225][6] ), .B2(n7495), 
        .Z(n1059) );
  OA22D0 U7051 ( .A1(n7496), .A2(prog_data[5]), .B1(\mem[225][5] ), .B2(n7495), 
        .Z(n1058) );
  OA22D0 U7052 ( .A1(n7496), .A2(prog_data[4]), .B1(\mem[225][4] ), .B2(n7495), 
        .Z(n1057) );
  OA22D0 U7053 ( .A1(n7496), .A2(prog_data[3]), .B1(\mem[225][3] ), .B2(n7495), 
        .Z(n1056) );
  OA22D0 U7054 ( .A1(n7496), .A2(prog_data[2]), .B1(\mem[225][2] ), .B2(n7495), 
        .Z(n1055) );
  OA22D0 U7055 ( .A1(n7496), .A2(prog_data[1]), .B1(\mem[225][1] ), .B2(n7495), 
        .Z(n1054) );
  OA22D0 U7056 ( .A1(n7496), .A2(prog_data[0]), .B1(\mem[225][0] ), .B2(n7495), 
        .Z(n1053) );
  INVD0 U7057 ( .I(n7497), .ZN(n7498) );
  OA22D0 U7058 ( .A1(n7498), .A2(prog_data[15]), .B1(\mem[226][15] ), .B2(
        n7497), .Z(n1052) );
  OA22D0 U7059 ( .A1(n7498), .A2(prog_data[14]), .B1(\mem[226][14] ), .B2(
        n7497), .Z(n1051) );
  OA22D0 U7060 ( .A1(n7498), .A2(prog_data[13]), .B1(\mem[226][13] ), .B2(
        n7497), .Z(n1050) );
  OA22D0 U7061 ( .A1(n7498), .A2(prog_data[12]), .B1(\mem[226][12] ), .B2(
        n7497), .Z(n1049) );
  OA22D0 U7062 ( .A1(n7498), .A2(prog_data[11]), .B1(\mem[226][11] ), .B2(
        n7497), .Z(n1048) );
  OA22D0 U7063 ( .A1(n7498), .A2(prog_data[10]), .B1(\mem[226][10] ), .B2(
        n7497), .Z(n1047) );
  OA22D0 U7064 ( .A1(n7498), .A2(prog_data[9]), .B1(\mem[226][9] ), .B2(n7497), 
        .Z(n1046) );
  OA22D0 U7065 ( .A1(n7498), .A2(prog_data[8]), .B1(\mem[226][8] ), .B2(n7497), 
        .Z(n1045) );
  OA22D0 U7066 ( .A1(n7498), .A2(prog_data[7]), .B1(\mem[226][7] ), .B2(n7497), 
        .Z(n1044) );
  OA22D0 U7067 ( .A1(n7498), .A2(prog_data[6]), .B1(\mem[226][6] ), .B2(n7497), 
        .Z(n1043) );
  OA22D0 U7068 ( .A1(n7498), .A2(prog_data[5]), .B1(\mem[226][5] ), .B2(n7497), 
        .Z(n1042) );
  OA22D0 U7069 ( .A1(n7498), .A2(prog_data[4]), .B1(\mem[226][4] ), .B2(n7497), 
        .Z(n1041) );
  OA22D0 U7070 ( .A1(n7498), .A2(prog_data[3]), .B1(\mem[226][3] ), .B2(n7497), 
        .Z(n1040) );
  OA22D0 U7071 ( .A1(n7498), .A2(prog_data[2]), .B1(\mem[226][2] ), .B2(n7497), 
        .Z(n1039) );
  OA22D0 U7072 ( .A1(n7498), .A2(prog_data[1]), .B1(\mem[226][1] ), .B2(n7497), 
        .Z(n1038) );
  OA22D0 U7073 ( .A1(n7498), .A2(prog_data[0]), .B1(\mem[226][0] ), .B2(n7497), 
        .Z(n1037) );
  NR2D0 U7074 ( .A1(n7537), .A2(n7523), .ZN(n7499) );
  INVD0 U7075 ( .I(n7499), .ZN(n7500) );
  OA22D0 U7076 ( .A1(n7500), .A2(prog_data[15]), .B1(\mem[227][15] ), .B2(
        n7499), .Z(n1036) );
  OA22D0 U7077 ( .A1(n7500), .A2(prog_data[14]), .B1(\mem[227][14] ), .B2(
        n7499), .Z(n1035) );
  OA22D0 U7078 ( .A1(n7500), .A2(prog_data[13]), .B1(\mem[227][13] ), .B2(
        n7499), .Z(n1034) );
  OA22D0 U7079 ( .A1(n7500), .A2(prog_data[12]), .B1(\mem[227][12] ), .B2(
        n7499), .Z(n1033) );
  OA22D0 U7080 ( .A1(n7500), .A2(prog_data[11]), .B1(\mem[227][11] ), .B2(
        n7499), .Z(n1032) );
  OA22D0 U7081 ( .A1(n7500), .A2(prog_data[10]), .B1(\mem[227][10] ), .B2(
        n7499), .Z(n1031) );
  OA22D0 U7082 ( .A1(n7500), .A2(prog_data[9]), .B1(\mem[227][9] ), .B2(n7499), 
        .Z(n1030) );
  OA22D0 U7083 ( .A1(n7500), .A2(prog_data[8]), .B1(\mem[227][8] ), .B2(n7499), 
        .Z(n1029) );
  OA22D0 U7084 ( .A1(n7500), .A2(prog_data[7]), .B1(\mem[227][7] ), .B2(n7499), 
        .Z(n1028) );
  OA22D0 U7085 ( .A1(n7500), .A2(prog_data[6]), .B1(\mem[227][6] ), .B2(n7499), 
        .Z(n1027) );
  OA22D0 U7086 ( .A1(n7500), .A2(prog_data[5]), .B1(\mem[227][5] ), .B2(n7499), 
        .Z(n1026) );
  OA22D0 U7087 ( .A1(n7500), .A2(prog_data[4]), .B1(\mem[227][4] ), .B2(n7499), 
        .Z(n1025) );
  OA22D0 U7088 ( .A1(n7500), .A2(prog_data[3]), .B1(\mem[227][3] ), .B2(n7499), 
        .Z(n1024) );
  OA22D0 U7089 ( .A1(n7500), .A2(prog_data[2]), .B1(\mem[227][2] ), .B2(n7499), 
        .Z(n1023) );
  OA22D0 U7090 ( .A1(n7500), .A2(prog_data[1]), .B1(\mem[227][1] ), .B2(n7499), 
        .Z(n1022) );
  OA22D0 U7091 ( .A1(n7500), .A2(prog_data[0]), .B1(\mem[227][0] ), .B2(n7499), 
        .Z(n1021) );
  NR2D0 U7092 ( .A1(n7540), .A2(n7523), .ZN(n7501) );
  INVD0 U7093 ( .I(n7501), .ZN(n7502) );
  OA22D0 U7094 ( .A1(n7502), .A2(prog_data[15]), .B1(\mem[228][15] ), .B2(
        n7501), .Z(n1020) );
  OA22D0 U7095 ( .A1(n7502), .A2(prog_data[14]), .B1(\mem[228][14] ), .B2(
        n7501), .Z(n1019) );
  OA22D0 U7096 ( .A1(n7502), .A2(prog_data[13]), .B1(\mem[228][13] ), .B2(
        n7501), .Z(n1018) );
  OA22D0 U7097 ( .A1(n7502), .A2(prog_data[12]), .B1(\mem[228][12] ), .B2(
        n7501), .Z(n1017) );
  OA22D0 U7098 ( .A1(n7502), .A2(prog_data[11]), .B1(\mem[228][11] ), .B2(
        n7501), .Z(n1016) );
  OA22D0 U7099 ( .A1(n7502), .A2(prog_data[10]), .B1(\mem[228][10] ), .B2(
        n7501), .Z(n1015) );
  OA22D0 U7100 ( .A1(n7502), .A2(prog_data[9]), .B1(\mem[228][9] ), .B2(n7501), 
        .Z(n1014) );
  OA22D0 U7101 ( .A1(n7502), .A2(prog_data[8]), .B1(\mem[228][8] ), .B2(n7501), 
        .Z(n1013) );
  OA22D0 U7102 ( .A1(n7502), .A2(prog_data[7]), .B1(\mem[228][7] ), .B2(n7501), 
        .Z(n1012) );
  OA22D0 U7103 ( .A1(n7502), .A2(prog_data[6]), .B1(\mem[228][6] ), .B2(n7501), 
        .Z(n1011) );
  OA22D0 U7104 ( .A1(n7502), .A2(prog_data[5]), .B1(\mem[228][5] ), .B2(n7501), 
        .Z(n1010) );
  OA22D0 U7105 ( .A1(n7502), .A2(prog_data[4]), .B1(\mem[228][4] ), .B2(n7501), 
        .Z(n1009) );
  OA22D0 U7106 ( .A1(n7502), .A2(prog_data[3]), .B1(\mem[228][3] ), .B2(n7501), 
        .Z(n1008) );
  OA22D0 U7107 ( .A1(n7502), .A2(prog_data[2]), .B1(\mem[228][2] ), .B2(n7501), 
        .Z(n1007) );
  OA22D0 U7108 ( .A1(n7502), .A2(prog_data[1]), .B1(\mem[228][1] ), .B2(n7501), 
        .Z(n1006) );
  OA22D0 U7109 ( .A1(n7502), .A2(prog_data[0]), .B1(\mem[228][0] ), .B2(n7501), 
        .Z(n1005) );
  NR2D0 U7110 ( .A1(n7543), .A2(n7523), .ZN(n7503) );
  INVD0 U7111 ( .I(n7503), .ZN(n7504) );
  OA22D0 U7112 ( .A1(n7504), .A2(prog_data[15]), .B1(\mem[229][15] ), .B2(
        n7503), .Z(n1004) );
  OA22D0 U7113 ( .A1(n7504), .A2(prog_data[14]), .B1(\mem[229][14] ), .B2(
        n7503), .Z(n1003) );
  OA22D0 U7114 ( .A1(n7504), .A2(prog_data[13]), .B1(\mem[229][13] ), .B2(
        n7503), .Z(n1002) );
  OA22D0 U7115 ( .A1(n7504), .A2(prog_data[12]), .B1(\mem[229][12] ), .B2(
        n7503), .Z(n1001) );
  OA22D0 U7116 ( .A1(n7504), .A2(prog_data[11]), .B1(\mem[229][11] ), .B2(
        n7503), .Z(n1000) );
  OA22D0 U7117 ( .A1(n7504), .A2(prog_data[10]), .B1(\mem[229][10] ), .B2(
        n7503), .Z(n999) );
  OA22D0 U7118 ( .A1(n7504), .A2(prog_data[9]), .B1(\mem[229][9] ), .B2(n7503), 
        .Z(n998) );
  OA22D0 U7119 ( .A1(n7504), .A2(prog_data[8]), .B1(\mem[229][8] ), .B2(n7503), 
        .Z(n997) );
  OA22D0 U7120 ( .A1(n7504), .A2(prog_data[7]), .B1(\mem[229][7] ), .B2(n7503), 
        .Z(n996) );
  OA22D0 U7121 ( .A1(n7504), .A2(prog_data[6]), .B1(\mem[229][6] ), .B2(n7503), 
        .Z(n995) );
  OA22D0 U7122 ( .A1(n7504), .A2(prog_data[5]), .B1(\mem[229][5] ), .B2(n7503), 
        .Z(n994) );
  OA22D0 U7123 ( .A1(n7504), .A2(prog_data[4]), .B1(\mem[229][4] ), .B2(n7503), 
        .Z(n993) );
  OA22D0 U7124 ( .A1(n7504), .A2(prog_data[3]), .B1(\mem[229][3] ), .B2(n7503), 
        .Z(n992) );
  OA22D0 U7125 ( .A1(n7504), .A2(prog_data[2]), .B1(\mem[229][2] ), .B2(n7503), 
        .Z(n991) );
  OA22D0 U7126 ( .A1(n7504), .A2(prog_data[1]), .B1(\mem[229][1] ), .B2(n7503), 
        .Z(n990) );
  OA22D0 U7127 ( .A1(n7504), .A2(prog_data[0]), .B1(\mem[229][0] ), .B2(n7503), 
        .Z(n989) );
  NR2D0 U7128 ( .A1(n7546), .A2(n7523), .ZN(n7505) );
  INVD0 U7129 ( .I(n7505), .ZN(n7506) );
  OA22D0 U7130 ( .A1(n7506), .A2(prog_data[15]), .B1(\mem[230][15] ), .B2(
        n7505), .Z(n988) );
  OA22D0 U7131 ( .A1(n7506), .A2(prog_data[14]), .B1(\mem[230][14] ), .B2(
        n7505), .Z(n987) );
  OA22D0 U7132 ( .A1(n7506), .A2(prog_data[13]), .B1(\mem[230][13] ), .B2(
        n7505), .Z(n986) );
  OA22D0 U7133 ( .A1(n7506), .A2(prog_data[12]), .B1(\mem[230][12] ), .B2(
        n7505), .Z(n985) );
  OA22D0 U7134 ( .A1(n7506), .A2(prog_data[11]), .B1(\mem[230][11] ), .B2(
        n7505), .Z(n984) );
  OA22D0 U7135 ( .A1(n7506), .A2(prog_data[10]), .B1(\mem[230][10] ), .B2(
        n7505), .Z(n983) );
  OA22D0 U7136 ( .A1(n7506), .A2(prog_data[9]), .B1(\mem[230][9] ), .B2(n7505), 
        .Z(n982) );
  OA22D0 U7137 ( .A1(n7506), .A2(prog_data[8]), .B1(\mem[230][8] ), .B2(n7505), 
        .Z(n981) );
  OA22D0 U7138 ( .A1(n7506), .A2(prog_data[7]), .B1(\mem[230][7] ), .B2(n7505), 
        .Z(n980) );
  OA22D0 U7139 ( .A1(n7506), .A2(prog_data[6]), .B1(\mem[230][6] ), .B2(n7505), 
        .Z(n979) );
  OA22D0 U7140 ( .A1(n7506), .A2(prog_data[5]), .B1(\mem[230][5] ), .B2(n7505), 
        .Z(n978) );
  OA22D0 U7141 ( .A1(n7506), .A2(prog_data[4]), .B1(\mem[230][4] ), .B2(n7505), 
        .Z(n977) );
  OA22D0 U7142 ( .A1(n7506), .A2(prog_data[3]), .B1(\mem[230][3] ), .B2(n7505), 
        .Z(n976) );
  OA22D0 U7143 ( .A1(n7506), .A2(prog_data[2]), .B1(\mem[230][2] ), .B2(n7505), 
        .Z(n975) );
  OA22D0 U7144 ( .A1(n7506), .A2(prog_data[1]), .B1(\mem[230][1] ), .B2(n7505), 
        .Z(n974) );
  OA22D0 U7145 ( .A1(n7506), .A2(prog_data[0]), .B1(\mem[230][0] ), .B2(n7505), 
        .Z(n973) );
  NR2D0 U7146 ( .A1(n7549), .A2(n7523), .ZN(n7507) );
  INVD0 U7147 ( .I(n7507), .ZN(n7508) );
  OA22D0 U7148 ( .A1(n7508), .A2(prog_data[15]), .B1(\mem[231][15] ), .B2(
        n7507), .Z(n972) );
  OA22D0 U7149 ( .A1(n7508), .A2(prog_data[14]), .B1(\mem[231][14] ), .B2(
        n7507), .Z(n971) );
  OA22D0 U7150 ( .A1(n7508), .A2(prog_data[13]), .B1(\mem[231][13] ), .B2(
        n7507), .Z(n970) );
  OA22D0 U7151 ( .A1(n7508), .A2(prog_data[12]), .B1(\mem[231][12] ), .B2(
        n7507), .Z(n969) );
  OA22D0 U7152 ( .A1(n7508), .A2(prog_data[11]), .B1(\mem[231][11] ), .B2(
        n7507), .Z(n968) );
  OA22D0 U7153 ( .A1(n7508), .A2(prog_data[10]), .B1(\mem[231][10] ), .B2(
        n7507), .Z(n967) );
  OA22D0 U7154 ( .A1(n7508), .A2(prog_data[9]), .B1(\mem[231][9] ), .B2(n7507), 
        .Z(n966) );
  OA22D0 U7155 ( .A1(n7508), .A2(prog_data[8]), .B1(\mem[231][8] ), .B2(n7507), 
        .Z(n965) );
  OA22D0 U7156 ( .A1(n7508), .A2(prog_data[7]), .B1(\mem[231][7] ), .B2(n7507), 
        .Z(n964) );
  OA22D0 U7157 ( .A1(n7508), .A2(prog_data[6]), .B1(\mem[231][6] ), .B2(n7507), 
        .Z(n963) );
  OA22D0 U7158 ( .A1(n7508), .A2(prog_data[5]), .B1(\mem[231][5] ), .B2(n7507), 
        .Z(n962) );
  OA22D0 U7159 ( .A1(n7508), .A2(prog_data[4]), .B1(\mem[231][4] ), .B2(n7507), 
        .Z(n961) );
  OA22D0 U7160 ( .A1(n7508), .A2(prog_data[3]), .B1(\mem[231][3] ), .B2(n7507), 
        .Z(n960) );
  OA22D0 U7161 ( .A1(n7508), .A2(prog_data[2]), .B1(\mem[231][2] ), .B2(n7507), 
        .Z(n959) );
  OA22D0 U7162 ( .A1(n7508), .A2(prog_data[1]), .B1(\mem[231][1] ), .B2(n7507), 
        .Z(n958) );
  OA22D0 U7163 ( .A1(n7508), .A2(prog_data[0]), .B1(\mem[231][0] ), .B2(n7507), 
        .Z(n957) );
  NR2D0 U7164 ( .A1(n7552), .A2(n7523), .ZN(n7509) );
  INVD0 U7165 ( .I(n7509), .ZN(n7510) );
  OA22D0 U7166 ( .A1(n7510), .A2(prog_data[15]), .B1(\mem[232][15] ), .B2(
        n7509), .Z(n956) );
  OA22D0 U7167 ( .A1(n7510), .A2(prog_data[14]), .B1(\mem[232][14] ), .B2(
        n7509), .Z(n955) );
  OA22D0 U7168 ( .A1(n7510), .A2(prog_data[13]), .B1(\mem[232][13] ), .B2(
        n7509), .Z(n954) );
  OA22D0 U7169 ( .A1(n7510), .A2(prog_data[12]), .B1(\mem[232][12] ), .B2(
        n7509), .Z(n953) );
  OA22D0 U7170 ( .A1(n7510), .A2(prog_data[11]), .B1(\mem[232][11] ), .B2(
        n7509), .Z(n952) );
  OA22D0 U7171 ( .A1(n7510), .A2(prog_data[10]), .B1(\mem[232][10] ), .B2(
        n7509), .Z(n951) );
  OA22D0 U7172 ( .A1(n7510), .A2(prog_data[9]), .B1(\mem[232][9] ), .B2(n7509), 
        .Z(n950) );
  OA22D0 U7173 ( .A1(n7510), .A2(prog_data[8]), .B1(\mem[232][8] ), .B2(n7509), 
        .Z(n949) );
  OA22D0 U7174 ( .A1(n7510), .A2(prog_data[7]), .B1(\mem[232][7] ), .B2(n7509), 
        .Z(n948) );
  OA22D0 U7175 ( .A1(n7510), .A2(prog_data[6]), .B1(\mem[232][6] ), .B2(n7509), 
        .Z(n947) );
  OA22D0 U7176 ( .A1(n7510), .A2(prog_data[5]), .B1(\mem[232][5] ), .B2(n7509), 
        .Z(n946) );
  OA22D0 U7177 ( .A1(n7510), .A2(prog_data[4]), .B1(\mem[232][4] ), .B2(n7509), 
        .Z(n945) );
  OA22D0 U7178 ( .A1(n7510), .A2(prog_data[3]), .B1(\mem[232][3] ), .B2(n7509), 
        .Z(n944) );
  OA22D0 U7179 ( .A1(n7510), .A2(prog_data[2]), .B1(\mem[232][2] ), .B2(n7509), 
        .Z(n943) );
  OA22D0 U7180 ( .A1(n7510), .A2(prog_data[1]), .B1(\mem[232][1] ), .B2(n7509), 
        .Z(n942) );
  OA22D0 U7181 ( .A1(n7510), .A2(prog_data[0]), .B1(\mem[232][0] ), .B2(n7509), 
        .Z(n941) );
  NR2D0 U7182 ( .A1(n7555), .A2(n7523), .ZN(n7511) );
  INVD0 U7183 ( .I(n7511), .ZN(n7512) );
  OA22D0 U7184 ( .A1(n7512), .A2(prog_data[15]), .B1(\mem[233][15] ), .B2(
        n7511), .Z(n940) );
  OA22D0 U7185 ( .A1(n7512), .A2(prog_data[14]), .B1(\mem[233][14] ), .B2(
        n7511), .Z(n939) );
  OA22D0 U7186 ( .A1(n7512), .A2(prog_data[13]), .B1(\mem[233][13] ), .B2(
        n7511), .Z(n938) );
  OA22D0 U7187 ( .A1(n7512), .A2(prog_data[12]), .B1(\mem[233][12] ), .B2(
        n7511), .Z(n937) );
  OA22D0 U7188 ( .A1(n7512), .A2(prog_data[11]), .B1(\mem[233][11] ), .B2(
        n7511), .Z(n936) );
  OA22D0 U7189 ( .A1(n7512), .A2(prog_data[10]), .B1(\mem[233][10] ), .B2(
        n7511), .Z(n935) );
  OA22D0 U7190 ( .A1(n7512), .A2(prog_data[9]), .B1(\mem[233][9] ), .B2(n7511), 
        .Z(n934) );
  OA22D0 U7191 ( .A1(n7512), .A2(prog_data[8]), .B1(\mem[233][8] ), .B2(n7511), 
        .Z(n933) );
  OA22D0 U7192 ( .A1(n7512), .A2(prog_data[7]), .B1(\mem[233][7] ), .B2(n7511), 
        .Z(n932) );
  OA22D0 U7193 ( .A1(n7512), .A2(prog_data[6]), .B1(\mem[233][6] ), .B2(n7511), 
        .Z(n931) );
  OA22D0 U7194 ( .A1(n7512), .A2(prog_data[5]), .B1(\mem[233][5] ), .B2(n7511), 
        .Z(n930) );
  OA22D0 U7195 ( .A1(n7512), .A2(prog_data[4]), .B1(\mem[233][4] ), .B2(n7511), 
        .Z(n929) );
  OA22D0 U7196 ( .A1(n7512), .A2(prog_data[3]), .B1(\mem[233][3] ), .B2(n7511), 
        .Z(n928) );
  OA22D0 U7197 ( .A1(n7512), .A2(prog_data[2]), .B1(\mem[233][2] ), .B2(n7511), 
        .Z(n927) );
  OA22D0 U7198 ( .A1(n7512), .A2(prog_data[1]), .B1(\mem[233][1] ), .B2(n7511), 
        .Z(n926) );
  OA22D0 U7199 ( .A1(n7512), .A2(prog_data[0]), .B1(\mem[233][0] ), .B2(n7511), 
        .Z(n925) );
  NR2D0 U7200 ( .A1(n7558), .A2(n7523), .ZN(n7513) );
  OA22D0 U7201 ( .A1(n7514), .A2(prog_data[15]), .B1(\mem[234][15] ), .B2(
        n7513), .Z(n924) );
  OA22D0 U7202 ( .A1(n7514), .A2(prog_data[14]), .B1(\mem[234][14] ), .B2(
        n7513), .Z(n923) );
  OA22D0 U7203 ( .A1(n7514), .A2(prog_data[13]), .B1(\mem[234][13] ), .B2(
        n7513), .Z(n922) );
  OA22D0 U7204 ( .A1(n7514), .A2(prog_data[12]), .B1(\mem[234][12] ), .B2(
        n7513), .Z(n921) );
  OA22D0 U7205 ( .A1(n7514), .A2(prog_data[11]), .B1(\mem[234][11] ), .B2(
        n7513), .Z(n920) );
  OA22D0 U7206 ( .A1(n7514), .A2(prog_data[10]), .B1(\mem[234][10] ), .B2(
        n7513), .Z(n919) );
  OA22D0 U7207 ( .A1(n7514), .A2(prog_data[9]), .B1(\mem[234][9] ), .B2(n7513), 
        .Z(n918) );
  OA22D0 U7208 ( .A1(n7514), .A2(prog_data[8]), .B1(\mem[234][8] ), .B2(n7513), 
        .Z(n917) );
  OA22D0 U7209 ( .A1(n7514), .A2(prog_data[7]), .B1(\mem[234][7] ), .B2(n7513), 
        .Z(n916) );
  OA22D0 U7210 ( .A1(n7514), .A2(prog_data[6]), .B1(\mem[234][6] ), .B2(n7513), 
        .Z(n915) );
  OA22D0 U7211 ( .A1(n7514), .A2(prog_data[5]), .B1(\mem[234][5] ), .B2(n7513), 
        .Z(n914) );
  OA22D0 U7212 ( .A1(n7514), .A2(prog_data[4]), .B1(\mem[234][4] ), .B2(n7513), 
        .Z(n913) );
  OA22D0 U7213 ( .A1(n7514), .A2(prog_data[3]), .B1(\mem[234][3] ), .B2(n7513), 
        .Z(n912) );
  OA22D0 U7214 ( .A1(n7514), .A2(prog_data[2]), .B1(\mem[234][2] ), .B2(n7513), 
        .Z(n911) );
  OA22D0 U7215 ( .A1(n7514), .A2(prog_data[1]), .B1(\mem[234][1] ), .B2(n7513), 
        .Z(n910) );
  OA22D0 U7216 ( .A1(n7514), .A2(prog_data[0]), .B1(\mem[234][0] ), .B2(n7513), 
        .Z(n909) );
  NR2D0 U7217 ( .A1(n7561), .A2(n7523), .ZN(n7515) );
  INVD0 U7218 ( .I(n7515), .ZN(n7516) );
  OA22D0 U7219 ( .A1(n7516), .A2(prog_data[15]), .B1(\mem[235][15] ), .B2(
        n7515), .Z(n908) );
  OA22D0 U7220 ( .A1(n7516), .A2(prog_data[14]), .B1(\mem[235][14] ), .B2(
        n7515), .Z(n907) );
  OA22D0 U7221 ( .A1(n7516), .A2(prog_data[13]), .B1(\mem[235][13] ), .B2(
        n7515), .Z(n906) );
  OA22D0 U7222 ( .A1(n7516), .A2(prog_data[12]), .B1(\mem[235][12] ), .B2(
        n7515), .Z(n905) );
  OA22D0 U7223 ( .A1(n7516), .A2(prog_data[11]), .B1(\mem[235][11] ), .B2(
        n7515), .Z(n904) );
  OA22D0 U7224 ( .A1(n7516), .A2(prog_data[10]), .B1(\mem[235][10] ), .B2(
        n7515), .Z(n903) );
  OA22D0 U7225 ( .A1(n7516), .A2(prog_data[9]), .B1(\mem[235][9] ), .B2(n7515), 
        .Z(n902) );
  OA22D0 U7226 ( .A1(n7516), .A2(prog_data[8]), .B1(\mem[235][8] ), .B2(n7515), 
        .Z(n901) );
  OA22D0 U7227 ( .A1(n7516), .A2(prog_data[7]), .B1(\mem[235][7] ), .B2(n7515), 
        .Z(n900) );
  OA22D0 U7228 ( .A1(n7516), .A2(prog_data[6]), .B1(\mem[235][6] ), .B2(n7515), 
        .Z(n899) );
  OA22D0 U7229 ( .A1(n7516), .A2(prog_data[5]), .B1(\mem[235][5] ), .B2(n7515), 
        .Z(n898) );
  OA22D0 U7230 ( .A1(n7516), .A2(prog_data[4]), .B1(\mem[235][4] ), .B2(n7515), 
        .Z(n897) );
  OA22D0 U7231 ( .A1(n7516), .A2(prog_data[3]), .B1(\mem[235][3] ), .B2(n7515), 
        .Z(n896) );
  OA22D0 U7232 ( .A1(n7516), .A2(prog_data[2]), .B1(\mem[235][2] ), .B2(n7515), 
        .Z(n895) );
  OA22D0 U7233 ( .A1(n7516), .A2(prog_data[1]), .B1(\mem[235][1] ), .B2(n7515), 
        .Z(n894) );
  OA22D0 U7234 ( .A1(n7516), .A2(prog_data[0]), .B1(\mem[235][0] ), .B2(n7515), 
        .Z(n893) );
  NR2D0 U7235 ( .A1(n7564), .A2(n7523), .ZN(n7517) );
  INVD0 U7236 ( .I(n7517), .ZN(n7518) );
  OA22D0 U7237 ( .A1(n7518), .A2(prog_data[15]), .B1(\mem[236][15] ), .B2(
        n7517), .Z(n892) );
  OA22D0 U7238 ( .A1(n7518), .A2(prog_data[14]), .B1(\mem[236][14] ), .B2(
        n7517), .Z(n891) );
  OA22D0 U7239 ( .A1(n7518), .A2(prog_data[13]), .B1(\mem[236][13] ), .B2(
        n7517), .Z(n890) );
  OA22D0 U7240 ( .A1(n7518), .A2(prog_data[12]), .B1(\mem[236][12] ), .B2(
        n7517), .Z(n889) );
  OA22D0 U7241 ( .A1(n7518), .A2(prog_data[11]), .B1(\mem[236][11] ), .B2(
        n7517), .Z(n888) );
  OA22D0 U7242 ( .A1(n7518), .A2(prog_data[10]), .B1(\mem[236][10] ), .B2(
        n7517), .Z(n887) );
  OA22D0 U7243 ( .A1(n7518), .A2(prog_data[9]), .B1(\mem[236][9] ), .B2(n7517), 
        .Z(n886) );
  OA22D0 U7244 ( .A1(n7518), .A2(prog_data[8]), .B1(\mem[236][8] ), .B2(n7517), 
        .Z(n885) );
  OA22D0 U7245 ( .A1(n7518), .A2(prog_data[7]), .B1(\mem[236][7] ), .B2(n7517), 
        .Z(n884) );
  OA22D0 U7246 ( .A1(n7518), .A2(prog_data[6]), .B1(\mem[236][6] ), .B2(n7517), 
        .Z(n883) );
  OA22D0 U7247 ( .A1(n7518), .A2(prog_data[5]), .B1(\mem[236][5] ), .B2(n7517), 
        .Z(n882) );
  OA22D0 U7248 ( .A1(n7518), .A2(prog_data[4]), .B1(\mem[236][4] ), .B2(n7517), 
        .Z(n881) );
  OA22D0 U7249 ( .A1(n7518), .A2(prog_data[3]), .B1(\mem[236][3] ), .B2(n7517), 
        .Z(n880) );
  OA22D0 U7250 ( .A1(n7518), .A2(prog_data[2]), .B1(\mem[236][2] ), .B2(n7517), 
        .Z(n879) );
  OA22D0 U7251 ( .A1(n7518), .A2(prog_data[1]), .B1(\mem[236][1] ), .B2(n7517), 
        .Z(n878) );
  OA22D0 U7252 ( .A1(n7518), .A2(prog_data[0]), .B1(\mem[236][0] ), .B2(n7517), 
        .Z(n877) );
  NR2D0 U7253 ( .A1(n7567), .A2(n7523), .ZN(n7519) );
  INVD0 U7254 ( .I(n7519), .ZN(n7520) );
  OA22D0 U7255 ( .A1(n7520), .A2(prog_data[15]), .B1(\mem[237][15] ), .B2(
        n7519), .Z(n876) );
  OA22D0 U7256 ( .A1(n7520), .A2(prog_data[14]), .B1(\mem[237][14] ), .B2(
        n7519), .Z(n875) );
  OA22D0 U7257 ( .A1(n7520), .A2(prog_data[13]), .B1(\mem[237][13] ), .B2(
        n7519), .Z(n874) );
  OA22D0 U7258 ( .A1(n7520), .A2(prog_data[12]), .B1(\mem[237][12] ), .B2(
        n7519), .Z(n873) );
  OA22D0 U7259 ( .A1(n7520), .A2(prog_data[11]), .B1(\mem[237][11] ), .B2(
        n7519), .Z(n872) );
  OA22D0 U7260 ( .A1(n7520), .A2(prog_data[10]), .B1(\mem[237][10] ), .B2(
        n7519), .Z(n871) );
  OA22D0 U7261 ( .A1(n7520), .A2(prog_data[9]), .B1(\mem[237][9] ), .B2(n7519), 
        .Z(n870) );
  OA22D0 U7262 ( .A1(n7520), .A2(prog_data[8]), .B1(\mem[237][8] ), .B2(n7519), 
        .Z(n869) );
  OA22D0 U7263 ( .A1(n7520), .A2(prog_data[7]), .B1(\mem[237][7] ), .B2(n7519), 
        .Z(n868) );
  OA22D0 U7264 ( .A1(n7520), .A2(prog_data[6]), .B1(\mem[237][6] ), .B2(n7519), 
        .Z(n867) );
  OA22D0 U7265 ( .A1(n7520), .A2(prog_data[5]), .B1(\mem[237][5] ), .B2(n7519), 
        .Z(n866) );
  OA22D0 U7266 ( .A1(n7520), .A2(prog_data[4]), .B1(\mem[237][4] ), .B2(n7519), 
        .Z(n865) );
  OA22D0 U7267 ( .A1(n7520), .A2(prog_data[3]), .B1(\mem[237][3] ), .B2(n7519), 
        .Z(n864) );
  OA22D0 U7268 ( .A1(n7520), .A2(prog_data[2]), .B1(\mem[237][2] ), .B2(n7519), 
        .Z(n863) );
  OA22D0 U7269 ( .A1(n7520), .A2(prog_data[1]), .B1(\mem[237][1] ), .B2(n7519), 
        .Z(n862) );
  OA22D0 U7270 ( .A1(n7520), .A2(prog_data[0]), .B1(\mem[237][0] ), .B2(n7519), 
        .Z(n861) );
  NR2D0 U7271 ( .A1(n7570), .A2(n7523), .ZN(n7521) );
  INVD0 U7272 ( .I(n7521), .ZN(n7522) );
  OA22D0 U7273 ( .A1(n7522), .A2(prog_data[15]), .B1(\mem[238][15] ), .B2(
        n7521), .Z(n860) );
  OA22D0 U7274 ( .A1(n7522), .A2(prog_data[14]), .B1(\mem[238][14] ), .B2(
        n7521), .Z(n859) );
  OA22D0 U7275 ( .A1(n7522), .A2(prog_data[13]), .B1(\mem[238][13] ), .B2(
        n7521), .Z(n858) );
  OA22D0 U7276 ( .A1(n7522), .A2(prog_data[12]), .B1(\mem[238][12] ), .B2(
        n7521), .Z(n857) );
  OA22D0 U7277 ( .A1(n7522), .A2(prog_data[11]), .B1(\mem[238][11] ), .B2(
        n7521), .Z(n856) );
  OA22D0 U7278 ( .A1(n7522), .A2(prog_data[10]), .B1(\mem[238][10] ), .B2(
        n7521), .Z(n855) );
  OA22D0 U7279 ( .A1(n7522), .A2(prog_data[9]), .B1(\mem[238][9] ), .B2(n7521), 
        .Z(n854) );
  OA22D0 U7280 ( .A1(n7522), .A2(prog_data[8]), .B1(\mem[238][8] ), .B2(n7521), 
        .Z(n853) );
  OA22D0 U7281 ( .A1(n7522), .A2(prog_data[7]), .B1(\mem[238][7] ), .B2(n7521), 
        .Z(n852) );
  OA22D0 U7282 ( .A1(n7522), .A2(prog_data[6]), .B1(\mem[238][6] ), .B2(n7521), 
        .Z(n851) );
  OA22D0 U7283 ( .A1(n7522), .A2(prog_data[5]), .B1(\mem[238][5] ), .B2(n7521), 
        .Z(n850) );
  OA22D0 U7284 ( .A1(n7522), .A2(prog_data[4]), .B1(\mem[238][4] ), .B2(n7521), 
        .Z(n849) );
  OA22D0 U7285 ( .A1(n7522), .A2(prog_data[3]), .B1(\mem[238][3] ), .B2(n7521), 
        .Z(n848) );
  OA22D0 U7286 ( .A1(n7522), .A2(prog_data[2]), .B1(\mem[238][2] ), .B2(n7521), 
        .Z(n847) );
  OA22D0 U7287 ( .A1(n7522), .A2(prog_data[1]), .B1(\mem[238][1] ), .B2(n7521), 
        .Z(n846) );
  OA22D0 U7288 ( .A1(n7522), .A2(prog_data[0]), .B1(\mem[238][0] ), .B2(n7521), 
        .Z(n845) );
  NR2D0 U7289 ( .A1(n7574), .A2(n7523), .ZN(n7524) );
  INVD0 U7290 ( .I(n7524), .ZN(n7525) );
  OA22D0 U7291 ( .A1(n7525), .A2(prog_data[15]), .B1(\mem[239][15] ), .B2(
        n7524), .Z(n844) );
  OA22D0 U7292 ( .A1(n7525), .A2(prog_data[14]), .B1(\mem[239][14] ), .B2(
        n7524), .Z(n843) );
  OA22D0 U7293 ( .A1(n7525), .A2(prog_data[13]), .B1(\mem[239][13] ), .B2(
        n7524), .Z(n842) );
  OA22D0 U7294 ( .A1(n7525), .A2(prog_data[12]), .B1(\mem[239][12] ), .B2(
        n7524), .Z(n841) );
  OA22D0 U7295 ( .A1(n7525), .A2(prog_data[11]), .B1(\mem[239][11] ), .B2(
        n7524), .Z(n840) );
  OA22D0 U7296 ( .A1(n7525), .A2(prog_data[10]), .B1(\mem[239][10] ), .B2(
        n7524), .Z(n839) );
  OA22D0 U7297 ( .A1(n7525), .A2(prog_data[9]), .B1(\mem[239][9] ), .B2(n7524), 
        .Z(n838) );
  OA22D0 U7298 ( .A1(n7525), .A2(prog_data[8]), .B1(\mem[239][8] ), .B2(n7524), 
        .Z(n837) );
  OA22D0 U7299 ( .A1(n7525), .A2(prog_data[7]), .B1(\mem[239][7] ), .B2(n7524), 
        .Z(n836) );
  OA22D0 U7300 ( .A1(n7525), .A2(prog_data[6]), .B1(\mem[239][6] ), .B2(n7524), 
        .Z(n835) );
  OA22D0 U7301 ( .A1(n7525), .A2(prog_data[5]), .B1(\mem[239][5] ), .B2(n7524), 
        .Z(n834) );
  OA22D0 U7302 ( .A1(n7525), .A2(prog_data[4]), .B1(\mem[239][4] ), .B2(n7524), 
        .Z(n833) );
  OA22D0 U7303 ( .A1(n7525), .A2(prog_data[3]), .B1(\mem[239][3] ), .B2(n7524), 
        .Z(n832) );
  OA22D0 U7304 ( .A1(n7525), .A2(prog_data[2]), .B1(\mem[239][2] ), .B2(n7524), 
        .Z(n831) );
  OA22D0 U7305 ( .A1(n7525), .A2(prog_data[1]), .B1(\mem[239][1] ), .B2(n7524), 
        .Z(n830) );
  OA22D0 U7306 ( .A1(n7525), .A2(prog_data[0]), .B1(\mem[239][0] ), .B2(n7524), 
        .Z(n829) );
  IND3D0 U7307 ( .A1(n7527), .B1(prog_addr[6]), .B2(n7526), .ZN(n7573) );
  NR2D0 U7308 ( .A1(n7528), .A2(n7573), .ZN(n7529) );
  INVD0 U7309 ( .I(n7529), .ZN(n7530) );
  OA22D0 U7310 ( .A1(n7530), .A2(prog_data[15]), .B1(\mem[240][15] ), .B2(
        n7529), .Z(n828) );
  OA22D0 U7311 ( .A1(n7530), .A2(prog_data[14]), .B1(\mem[240][14] ), .B2(
        n7529), .Z(n827) );
  OA22D0 U7312 ( .A1(n7530), .A2(prog_data[13]), .B1(\mem[240][13] ), .B2(
        n7529), .Z(n826) );
  OA22D0 U7313 ( .A1(n7530), .A2(prog_data[12]), .B1(\mem[240][12] ), .B2(
        n7529), .Z(n825) );
  OA22D0 U7314 ( .A1(n7530), .A2(prog_data[11]), .B1(\mem[240][11] ), .B2(
        n7529), .Z(n824) );
  OA22D0 U7315 ( .A1(n7530), .A2(prog_data[10]), .B1(\mem[240][10] ), .B2(
        n7529), .Z(n823) );
  OA22D0 U7316 ( .A1(n7530), .A2(prog_data[9]), .B1(\mem[240][9] ), .B2(n7529), 
        .Z(n822) );
  OA22D0 U7317 ( .A1(n7530), .A2(prog_data[8]), .B1(\mem[240][8] ), .B2(n7529), 
        .Z(n821) );
  OA22D0 U7318 ( .A1(n7530), .A2(prog_data[7]), .B1(\mem[240][7] ), .B2(n7529), 
        .Z(n820) );
  OA22D0 U7319 ( .A1(n7530), .A2(prog_data[6]), .B1(\mem[240][6] ), .B2(n7529), 
        .Z(n819) );
  OA22D0 U7320 ( .A1(n7530), .A2(prog_data[5]), .B1(\mem[240][5] ), .B2(n7529), 
        .Z(n818) );
  OA22D0 U7321 ( .A1(n7530), .A2(prog_data[4]), .B1(\mem[240][4] ), .B2(n7529), 
        .Z(n817) );
  OA22D0 U7322 ( .A1(n7530), .A2(prog_data[3]), .B1(\mem[240][3] ), .B2(n7529), 
        .Z(n816) );
  OA22D0 U7323 ( .A1(n7530), .A2(prog_data[2]), .B1(\mem[240][2] ), .B2(n7529), 
        .Z(n815) );
  OA22D0 U7324 ( .A1(n7530), .A2(prog_data[1]), .B1(\mem[240][1] ), .B2(n7529), 
        .Z(n814) );
  OA22D0 U7325 ( .A1(n7530), .A2(prog_data[0]), .B1(\mem[240][0] ), .B2(n7529), 
        .Z(n813) );
  INVD0 U7326 ( .I(n7532), .ZN(n7533) );
  OA22D0 U7327 ( .A1(n7533), .A2(prog_data[15]), .B1(\mem[241][15] ), .B2(
        n7532), .Z(n812) );
  OA22D0 U7328 ( .A1(n7533), .A2(prog_data[14]), .B1(\mem[241][14] ), .B2(
        n7532), .Z(n811) );
  OA22D0 U7329 ( .A1(n7533), .A2(prog_data[13]), .B1(\mem[241][13] ), .B2(
        n7532), .Z(n810) );
  OA22D0 U7330 ( .A1(n7533), .A2(prog_data[12]), .B1(\mem[241][12] ), .B2(
        n7532), .Z(n809) );
  OA22D0 U7331 ( .A1(n7533), .A2(prog_data[11]), .B1(\mem[241][11] ), .B2(
        n7532), .Z(n808) );
  OA22D0 U7332 ( .A1(n7533), .A2(prog_data[10]), .B1(\mem[241][10] ), .B2(
        n7532), .Z(n807) );
  OA22D0 U7333 ( .A1(n7533), .A2(prog_data[9]), .B1(\mem[241][9] ), .B2(n7532), 
        .Z(n806) );
  OA22D0 U7334 ( .A1(n7533), .A2(prog_data[8]), .B1(\mem[241][8] ), .B2(n7532), 
        .Z(n805) );
  OA22D0 U7335 ( .A1(n7533), .A2(prog_data[7]), .B1(\mem[241][7] ), .B2(n7532), 
        .Z(n804) );
  OA22D0 U7336 ( .A1(n7533), .A2(prog_data[6]), .B1(\mem[241][6] ), .B2(n7532), 
        .Z(n803) );
  OA22D0 U7337 ( .A1(n7533), .A2(prog_data[5]), .B1(\mem[241][5] ), .B2(n7532), 
        .Z(n802) );
  OA22D0 U7338 ( .A1(n7533), .A2(prog_data[4]), .B1(\mem[241][4] ), .B2(n7532), 
        .Z(n801) );
  OA22D0 U7339 ( .A1(n7533), .A2(prog_data[3]), .B1(\mem[241][3] ), .B2(n7532), 
        .Z(n800) );
  OA22D0 U7340 ( .A1(n7533), .A2(prog_data[2]), .B1(\mem[241][2] ), .B2(n7532), 
        .Z(n799) );
  OA22D0 U7341 ( .A1(n7533), .A2(prog_data[1]), .B1(\mem[241][1] ), .B2(n7532), 
        .Z(n798) );
  OA22D0 U7342 ( .A1(n7533), .A2(prog_data[0]), .B1(\mem[241][0] ), .B2(n7532), 
        .Z(n797) );
  NR2D0 U7343 ( .A1(n7534), .A2(n7573), .ZN(n7535) );
  INVD0 U7344 ( .I(n7535), .ZN(n7536) );
  OA22D0 U7345 ( .A1(n7536), .A2(prog_data[15]), .B1(\mem[242][15] ), .B2(
        n7535), .Z(n796) );
  OA22D0 U7346 ( .A1(n7536), .A2(prog_data[14]), .B1(\mem[242][14] ), .B2(
        n7535), .Z(n795) );
  OA22D0 U7347 ( .A1(n7536), .A2(prog_data[13]), .B1(\mem[242][13] ), .B2(
        n7535), .Z(n794) );
  OA22D0 U7348 ( .A1(n7536), .A2(prog_data[12]), .B1(\mem[242][12] ), .B2(
        n7535), .Z(n793) );
  OA22D0 U7349 ( .A1(n7536), .A2(prog_data[11]), .B1(\mem[242][11] ), .B2(
        n7535), .Z(n792) );
  OA22D0 U7350 ( .A1(n7536), .A2(prog_data[10]), .B1(\mem[242][10] ), .B2(
        n7535), .Z(n791) );
  OA22D0 U7351 ( .A1(n7536), .A2(prog_data[9]), .B1(\mem[242][9] ), .B2(n7535), 
        .Z(n790) );
  OA22D0 U7352 ( .A1(n7536), .A2(prog_data[8]), .B1(\mem[242][8] ), .B2(n7535), 
        .Z(n789) );
  OA22D0 U7353 ( .A1(n7536), .A2(prog_data[7]), .B1(\mem[242][7] ), .B2(n7535), 
        .Z(n788) );
  OA22D0 U7354 ( .A1(n7536), .A2(prog_data[6]), .B1(\mem[242][6] ), .B2(n7535), 
        .Z(n787) );
  OA22D0 U7355 ( .A1(n7536), .A2(prog_data[5]), .B1(\mem[242][5] ), .B2(n7535), 
        .Z(n786) );
  OA22D0 U7356 ( .A1(n7536), .A2(prog_data[4]), .B1(\mem[242][4] ), .B2(n7535), 
        .Z(n785) );
  OA22D0 U7357 ( .A1(n7536), .A2(prog_data[3]), .B1(\mem[242][3] ), .B2(n7535), 
        .Z(n784) );
  OA22D0 U7358 ( .A1(n7536), .A2(prog_data[2]), .B1(\mem[242][2] ), .B2(n7535), 
        .Z(n783) );
  OA22D0 U7359 ( .A1(n7536), .A2(prog_data[1]), .B1(\mem[242][1] ), .B2(n7535), 
        .Z(n782) );
  OA22D0 U7360 ( .A1(n7536), .A2(prog_data[0]), .B1(\mem[242][0] ), .B2(n7535), 
        .Z(n781) );
  NR2D0 U7361 ( .A1(n7537), .A2(n7573), .ZN(n7538) );
  INVD0 U7362 ( .I(n7538), .ZN(n7539) );
  OA22D0 U7363 ( .A1(n7539), .A2(prog_data[15]), .B1(\mem[243][15] ), .B2(
        n7538), .Z(n780) );
  OA22D0 U7364 ( .A1(n7539), .A2(prog_data[14]), .B1(\mem[243][14] ), .B2(
        n7538), .Z(n779) );
  OA22D0 U7365 ( .A1(n7539), .A2(prog_data[13]), .B1(\mem[243][13] ), .B2(
        n7538), .Z(n778) );
  OA22D0 U7366 ( .A1(n7539), .A2(prog_data[12]), .B1(\mem[243][12] ), .B2(
        n7538), .Z(n777) );
  OA22D0 U7367 ( .A1(n7539), .A2(prog_data[11]), .B1(\mem[243][11] ), .B2(
        n7538), .Z(n776) );
  OA22D0 U7368 ( .A1(n7539), .A2(prog_data[10]), .B1(\mem[243][10] ), .B2(
        n7538), .Z(n775) );
  OA22D0 U7369 ( .A1(n7539), .A2(prog_data[9]), .B1(\mem[243][9] ), .B2(n7538), 
        .Z(n774) );
  OA22D0 U7370 ( .A1(n7539), .A2(prog_data[8]), .B1(\mem[243][8] ), .B2(n7538), 
        .Z(n773) );
  OA22D0 U7371 ( .A1(n7539), .A2(prog_data[7]), .B1(\mem[243][7] ), .B2(n7538), 
        .Z(n772) );
  OA22D0 U7372 ( .A1(n7539), .A2(prog_data[6]), .B1(\mem[243][6] ), .B2(n7538), 
        .Z(n771) );
  OA22D0 U7373 ( .A1(n7539), .A2(prog_data[5]), .B1(\mem[243][5] ), .B2(n7538), 
        .Z(n770) );
  OA22D0 U7374 ( .A1(n7539), .A2(prog_data[4]), .B1(\mem[243][4] ), .B2(n7538), 
        .Z(n769) );
  OA22D0 U7375 ( .A1(n7539), .A2(prog_data[3]), .B1(\mem[243][3] ), .B2(n7538), 
        .Z(n768) );
  OA22D0 U7376 ( .A1(n7539), .A2(prog_data[2]), .B1(\mem[243][2] ), .B2(n7538), 
        .Z(n767) );
  OA22D0 U7377 ( .A1(n7539), .A2(prog_data[1]), .B1(\mem[243][1] ), .B2(n7538), 
        .Z(n766) );
  OA22D0 U7378 ( .A1(n7539), .A2(prog_data[0]), .B1(\mem[243][0] ), .B2(n7538), 
        .Z(n765) );
  NR2D0 U7379 ( .A1(n7540), .A2(n7573), .ZN(n7541) );
  INVD0 U7380 ( .I(n7541), .ZN(n7542) );
  OA22D0 U7381 ( .A1(n7542), .A2(prog_data[15]), .B1(\mem[244][15] ), .B2(
        n7541), .Z(n764) );
  OA22D0 U7382 ( .A1(n7542), .A2(prog_data[14]), .B1(\mem[244][14] ), .B2(
        n7541), .Z(n763) );
  OA22D0 U7383 ( .A1(n7542), .A2(prog_data[13]), .B1(\mem[244][13] ), .B2(
        n7541), .Z(n762) );
  OA22D0 U7384 ( .A1(n7542), .A2(prog_data[12]), .B1(\mem[244][12] ), .B2(
        n7541), .Z(n761) );
  OA22D0 U7385 ( .A1(n7542), .A2(prog_data[11]), .B1(\mem[244][11] ), .B2(
        n7541), .Z(n760) );
  OA22D0 U7386 ( .A1(n7542), .A2(prog_data[10]), .B1(\mem[244][10] ), .B2(
        n7541), .Z(n759) );
  OA22D0 U7387 ( .A1(n7542), .A2(prog_data[9]), .B1(\mem[244][9] ), .B2(n7541), 
        .Z(n758) );
  OA22D0 U7388 ( .A1(n7542), .A2(prog_data[8]), .B1(\mem[244][8] ), .B2(n7541), 
        .Z(n757) );
  OA22D0 U7389 ( .A1(n7542), .A2(prog_data[7]), .B1(\mem[244][7] ), .B2(n7541), 
        .Z(n756) );
  OA22D0 U7390 ( .A1(n7542), .A2(prog_data[6]), .B1(\mem[244][6] ), .B2(n7541), 
        .Z(n755) );
  OA22D0 U7391 ( .A1(n7542), .A2(prog_data[5]), .B1(\mem[244][5] ), .B2(n7541), 
        .Z(n754) );
  OA22D0 U7392 ( .A1(n7542), .A2(prog_data[4]), .B1(\mem[244][4] ), .B2(n7541), 
        .Z(n753) );
  OA22D0 U7393 ( .A1(n7542), .A2(prog_data[3]), .B1(\mem[244][3] ), .B2(n7541), 
        .Z(n752) );
  OA22D0 U7394 ( .A1(n7542), .A2(prog_data[2]), .B1(\mem[244][2] ), .B2(n7541), 
        .Z(n751) );
  OA22D0 U7395 ( .A1(n7542), .A2(prog_data[1]), .B1(\mem[244][1] ), .B2(n7541), 
        .Z(n750) );
  OA22D0 U7396 ( .A1(n7542), .A2(prog_data[0]), .B1(\mem[244][0] ), .B2(n7541), 
        .Z(n749) );
  NR2D0 U7397 ( .A1(n7543), .A2(n7573), .ZN(n7544) );
  INVD0 U7398 ( .I(n7544), .ZN(n7545) );
  OA22D0 U7399 ( .A1(n7545), .A2(prog_data[15]), .B1(\mem[245][15] ), .B2(
        n7544), .Z(n748) );
  OA22D0 U7400 ( .A1(n7545), .A2(prog_data[14]), .B1(\mem[245][14] ), .B2(
        n7544), .Z(n747) );
  OA22D0 U7401 ( .A1(n7545), .A2(prog_data[13]), .B1(\mem[245][13] ), .B2(
        n7544), .Z(n746) );
  OA22D0 U7402 ( .A1(n7545), .A2(prog_data[12]), .B1(\mem[245][12] ), .B2(
        n7544), .Z(n745) );
  OA22D0 U7403 ( .A1(n7545), .A2(prog_data[11]), .B1(\mem[245][11] ), .B2(
        n7544), .Z(n744) );
  OA22D0 U7404 ( .A1(n7545), .A2(prog_data[10]), .B1(\mem[245][10] ), .B2(
        n7544), .Z(n743) );
  OA22D0 U7405 ( .A1(n7545), .A2(prog_data[9]), .B1(\mem[245][9] ), .B2(n7544), 
        .Z(n742) );
  OA22D0 U7406 ( .A1(n7545), .A2(prog_data[8]), .B1(\mem[245][8] ), .B2(n7544), 
        .Z(n741) );
  OA22D0 U7407 ( .A1(n7545), .A2(prog_data[7]), .B1(\mem[245][7] ), .B2(n7544), 
        .Z(n740) );
  OA22D0 U7408 ( .A1(n7545), .A2(prog_data[6]), .B1(\mem[245][6] ), .B2(n7544), 
        .Z(n739) );
  OA22D0 U7409 ( .A1(n7545), .A2(prog_data[5]), .B1(\mem[245][5] ), .B2(n7544), 
        .Z(n738) );
  OA22D0 U7410 ( .A1(n7545), .A2(prog_data[4]), .B1(\mem[245][4] ), .B2(n7544), 
        .Z(n737) );
  OA22D0 U7411 ( .A1(n7545), .A2(prog_data[3]), .B1(\mem[245][3] ), .B2(n7544), 
        .Z(n736) );
  OA22D0 U7412 ( .A1(n7545), .A2(prog_data[2]), .B1(\mem[245][2] ), .B2(n7544), 
        .Z(n735) );
  OA22D0 U7413 ( .A1(n7545), .A2(prog_data[1]), .B1(\mem[245][1] ), .B2(n7544), 
        .Z(n734) );
  OA22D0 U7414 ( .A1(n7545), .A2(prog_data[0]), .B1(\mem[245][0] ), .B2(n7544), 
        .Z(n733) );
  NR2D0 U7415 ( .A1(n7546), .A2(n7573), .ZN(n7547) );
  INVD0 U7416 ( .I(n7547), .ZN(n7548) );
  OA22D0 U7417 ( .A1(n7548), .A2(prog_data[15]), .B1(\mem[246][15] ), .B2(
        n7547), .Z(n732) );
  OA22D0 U7418 ( .A1(n7548), .A2(prog_data[14]), .B1(\mem[246][14] ), .B2(
        n7547), .Z(n731) );
  OA22D0 U7419 ( .A1(n7548), .A2(prog_data[13]), .B1(\mem[246][13] ), .B2(
        n7547), .Z(n730) );
  OA22D0 U7420 ( .A1(n7548), .A2(prog_data[12]), .B1(\mem[246][12] ), .B2(
        n7547), .Z(n729) );
  OA22D0 U7421 ( .A1(n7548), .A2(prog_data[11]), .B1(\mem[246][11] ), .B2(
        n7547), .Z(n728) );
  OA22D0 U7422 ( .A1(n7548), .A2(prog_data[10]), .B1(\mem[246][10] ), .B2(
        n7547), .Z(n727) );
  OA22D0 U7423 ( .A1(n7548), .A2(prog_data[9]), .B1(\mem[246][9] ), .B2(n7547), 
        .Z(n726) );
  OA22D0 U7424 ( .A1(n7548), .A2(prog_data[8]), .B1(\mem[246][8] ), .B2(n7547), 
        .Z(n725) );
  OA22D0 U7425 ( .A1(n7548), .A2(prog_data[7]), .B1(\mem[246][7] ), .B2(n7547), 
        .Z(n724) );
  OA22D0 U7426 ( .A1(n7548), .A2(prog_data[6]), .B1(\mem[246][6] ), .B2(n7547), 
        .Z(n723) );
  OA22D0 U7427 ( .A1(n7548), .A2(prog_data[5]), .B1(\mem[246][5] ), .B2(n7547), 
        .Z(n722) );
  OA22D0 U7428 ( .A1(n7548), .A2(prog_data[4]), .B1(\mem[246][4] ), .B2(n7547), 
        .Z(n721) );
  OA22D0 U7429 ( .A1(n7548), .A2(prog_data[3]), .B1(\mem[246][3] ), .B2(n7547), 
        .Z(n720) );
  OA22D0 U7430 ( .A1(n7548), .A2(prog_data[2]), .B1(\mem[246][2] ), .B2(n7547), 
        .Z(n719) );
  OA22D0 U7431 ( .A1(n7548), .A2(prog_data[1]), .B1(\mem[246][1] ), .B2(n7547), 
        .Z(n718) );
  OA22D0 U7432 ( .A1(n7548), .A2(prog_data[0]), .B1(\mem[246][0] ), .B2(n7547), 
        .Z(n717) );
  NR2D0 U7433 ( .A1(n7549), .A2(n7573), .ZN(n7550) );
  INVD0 U7434 ( .I(n7550), .ZN(n7551) );
  OA22D0 U7435 ( .A1(n7551), .A2(prog_data[15]), .B1(\mem[247][15] ), .B2(
        n7550), .Z(n716) );
  OA22D0 U7436 ( .A1(n7551), .A2(prog_data[14]), .B1(\mem[247][14] ), .B2(
        n7550), .Z(n715) );
  OA22D0 U7437 ( .A1(n7551), .A2(prog_data[13]), .B1(\mem[247][13] ), .B2(
        n7550), .Z(n714) );
  OA22D0 U7438 ( .A1(n7551), .A2(prog_data[12]), .B1(\mem[247][12] ), .B2(
        n7550), .Z(n713) );
  OA22D0 U7439 ( .A1(n7551), .A2(prog_data[11]), .B1(\mem[247][11] ), .B2(
        n7550), .Z(n712) );
  OA22D0 U7440 ( .A1(n7551), .A2(prog_data[10]), .B1(\mem[247][10] ), .B2(
        n7550), .Z(n711) );
  OA22D0 U7441 ( .A1(n7551), .A2(prog_data[9]), .B1(\mem[247][9] ), .B2(n7550), 
        .Z(n710) );
  OA22D0 U7442 ( .A1(n7551), .A2(prog_data[8]), .B1(\mem[247][8] ), .B2(n7550), 
        .Z(n709) );
  OA22D0 U7443 ( .A1(n7551), .A2(prog_data[7]), .B1(\mem[247][7] ), .B2(n7550), 
        .Z(n708) );
  OA22D0 U7444 ( .A1(n7551), .A2(prog_data[6]), .B1(\mem[247][6] ), .B2(n7550), 
        .Z(n707) );
  OA22D0 U7445 ( .A1(n7551), .A2(prog_data[5]), .B1(\mem[247][5] ), .B2(n7550), 
        .Z(n706) );
  OA22D0 U7446 ( .A1(n7551), .A2(prog_data[4]), .B1(\mem[247][4] ), .B2(n7550), 
        .Z(n705) );
  OA22D0 U7447 ( .A1(n7551), .A2(prog_data[3]), .B1(\mem[247][3] ), .B2(n7550), 
        .Z(n704) );
  OA22D0 U7448 ( .A1(n7551), .A2(prog_data[2]), .B1(\mem[247][2] ), .B2(n7550), 
        .Z(n703) );
  OA22D0 U7449 ( .A1(n7551), .A2(prog_data[1]), .B1(\mem[247][1] ), .B2(n7550), 
        .Z(n702) );
  OA22D0 U7450 ( .A1(n7551), .A2(prog_data[0]), .B1(\mem[247][0] ), .B2(n7550), 
        .Z(n701) );
  NR2D0 U7451 ( .A1(n7552), .A2(n7573), .ZN(n7553) );
  INVD0 U7452 ( .I(n7553), .ZN(n7554) );
  OA22D0 U7453 ( .A1(n7554), .A2(prog_data[15]), .B1(\mem[248][15] ), .B2(
        n7553), .Z(n700) );
  OA22D0 U7454 ( .A1(n7554), .A2(prog_data[14]), .B1(\mem[248][14] ), .B2(
        n7553), .Z(n699) );
  OA22D0 U7455 ( .A1(n7554), .A2(prog_data[13]), .B1(\mem[248][13] ), .B2(
        n7553), .Z(n698) );
  OA22D0 U7456 ( .A1(n7554), .A2(prog_data[12]), .B1(\mem[248][12] ), .B2(
        n7553), .Z(n697) );
  OA22D0 U7457 ( .A1(n7554), .A2(prog_data[11]), .B1(\mem[248][11] ), .B2(
        n7553), .Z(n696) );
  OA22D0 U7458 ( .A1(n7554), .A2(prog_data[10]), .B1(\mem[248][10] ), .B2(
        n7553), .Z(n695) );
  OA22D0 U7459 ( .A1(n7554), .A2(prog_data[9]), .B1(\mem[248][9] ), .B2(n7553), 
        .Z(n694) );
  OA22D0 U7460 ( .A1(n7554), .A2(prog_data[8]), .B1(\mem[248][8] ), .B2(n7553), 
        .Z(n693) );
  OA22D0 U7461 ( .A1(n7554), .A2(prog_data[7]), .B1(\mem[248][7] ), .B2(n7553), 
        .Z(n692) );
  OA22D0 U7462 ( .A1(n7554), .A2(prog_data[6]), .B1(\mem[248][6] ), .B2(n7553), 
        .Z(n691) );
  OA22D0 U7463 ( .A1(n7554), .A2(prog_data[5]), .B1(\mem[248][5] ), .B2(n7553), 
        .Z(n690) );
  OA22D0 U7464 ( .A1(n7554), .A2(prog_data[4]), .B1(\mem[248][4] ), .B2(n7553), 
        .Z(n689) );
  OA22D0 U7465 ( .A1(n7554), .A2(prog_data[3]), .B1(\mem[248][3] ), .B2(n7553), 
        .Z(n688) );
  OA22D0 U7466 ( .A1(n7554), .A2(prog_data[2]), .B1(\mem[248][2] ), .B2(n7553), 
        .Z(n687) );
  OA22D0 U7467 ( .A1(n7554), .A2(prog_data[1]), .B1(\mem[248][1] ), .B2(n7553), 
        .Z(n686) );
  OA22D0 U7468 ( .A1(n7554), .A2(prog_data[0]), .B1(\mem[248][0] ), .B2(n7553), 
        .Z(n685) );
  NR2D0 U7469 ( .A1(n7555), .A2(n7573), .ZN(n7556) );
  OA22D0 U7470 ( .A1(n7557), .A2(prog_data[15]), .B1(\mem[249][15] ), .B2(
        n7556), .Z(n684) );
  OA22D0 U7471 ( .A1(n7557), .A2(prog_data[14]), .B1(\mem[249][14] ), .B2(
        n7556), .Z(n683) );
  OA22D0 U7472 ( .A1(n7557), .A2(prog_data[13]), .B1(\mem[249][13] ), .B2(
        n7556), .Z(n682) );
  OA22D0 U7473 ( .A1(n7557), .A2(prog_data[12]), .B1(\mem[249][12] ), .B2(
        n7556), .Z(n681) );
  OA22D0 U7474 ( .A1(n7557), .A2(prog_data[11]), .B1(\mem[249][11] ), .B2(
        n7556), .Z(n680) );
  OA22D0 U7475 ( .A1(n7557), .A2(prog_data[10]), .B1(\mem[249][10] ), .B2(
        n7556), .Z(n679) );
  OA22D0 U7476 ( .A1(n7557), .A2(prog_data[9]), .B1(\mem[249][9] ), .B2(n7556), 
        .Z(n678) );
  OA22D0 U7477 ( .A1(n7557), .A2(prog_data[8]), .B1(\mem[249][8] ), .B2(n7556), 
        .Z(n677) );
  OA22D0 U7478 ( .A1(n7557), .A2(prog_data[7]), .B1(\mem[249][7] ), .B2(n7556), 
        .Z(n676) );
  OA22D0 U7479 ( .A1(n7557), .A2(prog_data[6]), .B1(\mem[249][6] ), .B2(n7556), 
        .Z(n675) );
  OA22D0 U7480 ( .A1(n7557), .A2(prog_data[5]), .B1(\mem[249][5] ), .B2(n7556), 
        .Z(n674) );
  OA22D0 U7481 ( .A1(n7557), .A2(prog_data[4]), .B1(\mem[249][4] ), .B2(n7556), 
        .Z(n673) );
  OA22D0 U7482 ( .A1(n7557), .A2(prog_data[3]), .B1(\mem[249][3] ), .B2(n7556), 
        .Z(n672) );
  OA22D0 U7483 ( .A1(n7557), .A2(prog_data[2]), .B1(\mem[249][2] ), .B2(n7556), 
        .Z(n671) );
  OA22D0 U7484 ( .A1(n7557), .A2(prog_data[1]), .B1(\mem[249][1] ), .B2(n7556), 
        .Z(n670) );
  OA22D0 U7485 ( .A1(n7557), .A2(prog_data[0]), .B1(\mem[249][0] ), .B2(n7556), 
        .Z(n669) );
  NR2D0 U7486 ( .A1(n7558), .A2(n7573), .ZN(n7559) );
  INVD0 U7487 ( .I(n7559), .ZN(n7560) );
  OA22D0 U7488 ( .A1(n7560), .A2(prog_data[15]), .B1(\mem[250][15] ), .B2(
        n7559), .Z(n668) );
  OA22D0 U7489 ( .A1(n7560), .A2(prog_data[14]), .B1(\mem[250][14] ), .B2(
        n7559), .Z(n667) );
  OA22D0 U7490 ( .A1(n7560), .A2(prog_data[13]), .B1(\mem[250][13] ), .B2(
        n7559), .Z(n666) );
  OA22D0 U7491 ( .A1(n7560), .A2(prog_data[12]), .B1(\mem[250][12] ), .B2(
        n7559), .Z(n665) );
  OA22D0 U7492 ( .A1(n7560), .A2(prog_data[11]), .B1(\mem[250][11] ), .B2(
        n7559), .Z(n664) );
  OA22D0 U7493 ( .A1(n7560), .A2(prog_data[10]), .B1(\mem[250][10] ), .B2(
        n7559), .Z(n663) );
  OA22D0 U7494 ( .A1(n7560), .A2(prog_data[9]), .B1(\mem[250][9] ), .B2(n7559), 
        .Z(n662) );
  OA22D0 U7495 ( .A1(n7560), .A2(prog_data[8]), .B1(\mem[250][8] ), .B2(n7559), 
        .Z(n661) );
  OA22D0 U7496 ( .A1(n7560), .A2(prog_data[7]), .B1(\mem[250][7] ), .B2(n7559), 
        .Z(n660) );
  OA22D0 U7497 ( .A1(n7560), .A2(prog_data[6]), .B1(\mem[250][6] ), .B2(n7559), 
        .Z(n659) );
  OA22D0 U7498 ( .A1(n7560), .A2(prog_data[5]), .B1(\mem[250][5] ), .B2(n7559), 
        .Z(n658) );
  OA22D0 U7499 ( .A1(n7560), .A2(prog_data[4]), .B1(\mem[250][4] ), .B2(n7559), 
        .Z(n657) );
  OA22D0 U7500 ( .A1(n7560), .A2(prog_data[3]), .B1(\mem[250][3] ), .B2(n7559), 
        .Z(n656) );
  OA22D0 U7501 ( .A1(n7560), .A2(prog_data[2]), .B1(\mem[250][2] ), .B2(n7559), 
        .Z(n655) );
  OA22D0 U7502 ( .A1(n7560), .A2(prog_data[1]), .B1(\mem[250][1] ), .B2(n7559), 
        .Z(n654) );
  OA22D0 U7503 ( .A1(n7560), .A2(prog_data[0]), .B1(\mem[250][0] ), .B2(n7559), 
        .Z(n653) );
  NR2D0 U7504 ( .A1(n7561), .A2(n7573), .ZN(n7562) );
  INVD0 U7505 ( .I(n7562), .ZN(n7563) );
  OA22D0 U7506 ( .A1(n7563), .A2(prog_data[15]), .B1(\mem[251][15] ), .B2(
        n7562), .Z(n652) );
  OA22D0 U7507 ( .A1(n7563), .A2(prog_data[14]), .B1(\mem[251][14] ), .B2(
        n7562), .Z(n651) );
  OA22D0 U7508 ( .A1(n7563), .A2(prog_data[13]), .B1(\mem[251][13] ), .B2(
        n7562), .Z(n650) );
  OA22D0 U7509 ( .A1(n7563), .A2(prog_data[12]), .B1(\mem[251][12] ), .B2(
        n7562), .Z(n649) );
  OA22D0 U7510 ( .A1(n7563), .A2(prog_data[11]), .B1(\mem[251][11] ), .B2(
        n7562), .Z(n648) );
  OA22D0 U7511 ( .A1(n7563), .A2(prog_data[10]), .B1(\mem[251][10] ), .B2(
        n7562), .Z(n647) );
  OA22D0 U7512 ( .A1(n7563), .A2(prog_data[9]), .B1(\mem[251][9] ), .B2(n7562), 
        .Z(n646) );
  OA22D0 U7513 ( .A1(n7563), .A2(prog_data[8]), .B1(\mem[251][8] ), .B2(n7562), 
        .Z(n645) );
  OA22D0 U7514 ( .A1(n7563), .A2(prog_data[7]), .B1(\mem[251][7] ), .B2(n7562), 
        .Z(n644) );
  OA22D0 U7515 ( .A1(n7563), .A2(prog_data[6]), .B1(\mem[251][6] ), .B2(n7562), 
        .Z(n643) );
  OA22D0 U7516 ( .A1(n7563), .A2(prog_data[5]), .B1(\mem[251][5] ), .B2(n7562), 
        .Z(n642) );
  OA22D0 U7517 ( .A1(n7563), .A2(prog_data[4]), .B1(\mem[251][4] ), .B2(n7562), 
        .Z(n641) );
  OA22D0 U7518 ( .A1(n7563), .A2(prog_data[3]), .B1(\mem[251][3] ), .B2(n7562), 
        .Z(n640) );
  OA22D0 U7519 ( .A1(n7563), .A2(prog_data[2]), .B1(\mem[251][2] ), .B2(n7562), 
        .Z(n639) );
  OA22D0 U7520 ( .A1(n7563), .A2(prog_data[1]), .B1(\mem[251][1] ), .B2(n7562), 
        .Z(n638) );
  OA22D0 U7521 ( .A1(n7563), .A2(prog_data[0]), .B1(\mem[251][0] ), .B2(n7562), 
        .Z(n637) );
  NR2D0 U7522 ( .A1(n7564), .A2(n7573), .ZN(n7565) );
  INVD0 U7523 ( .I(n7565), .ZN(n7566) );
  OA22D0 U7524 ( .A1(n7566), .A2(prog_data[15]), .B1(\mem[252][15] ), .B2(
        n7565), .Z(n636) );
  OA22D0 U7525 ( .A1(n7566), .A2(prog_data[14]), .B1(\mem[252][14] ), .B2(
        n7565), .Z(n635) );
  OA22D0 U7526 ( .A1(n7566), .A2(prog_data[13]), .B1(\mem[252][13] ), .B2(
        n7565), .Z(n634) );
  OA22D0 U7527 ( .A1(n7566), .A2(prog_data[12]), .B1(\mem[252][12] ), .B2(
        n7565), .Z(n633) );
  OA22D0 U7528 ( .A1(n7566), .A2(prog_data[11]), .B1(\mem[252][11] ), .B2(
        n7565), .Z(n632) );
  OA22D0 U7529 ( .A1(n7566), .A2(prog_data[10]), .B1(\mem[252][10] ), .B2(
        n7565), .Z(n631) );
  OA22D0 U7530 ( .A1(n7566), .A2(prog_data[9]), .B1(\mem[252][9] ), .B2(n7565), 
        .Z(n630) );
  OA22D0 U7531 ( .A1(n7566), .A2(prog_data[8]), .B1(\mem[252][8] ), .B2(n7565), 
        .Z(n629) );
  OA22D0 U7532 ( .A1(n7566), .A2(prog_data[7]), .B1(\mem[252][7] ), .B2(n7565), 
        .Z(n628) );
  OA22D0 U7533 ( .A1(n7566), .A2(prog_data[6]), .B1(\mem[252][6] ), .B2(n7565), 
        .Z(n627) );
  OA22D0 U7534 ( .A1(n7566), .A2(prog_data[5]), .B1(\mem[252][5] ), .B2(n7565), 
        .Z(n626) );
  OA22D0 U7535 ( .A1(n7566), .A2(prog_data[4]), .B1(\mem[252][4] ), .B2(n7565), 
        .Z(n625) );
  OA22D0 U7536 ( .A1(n7566), .A2(prog_data[3]), .B1(\mem[252][3] ), .B2(n7565), 
        .Z(n624) );
  OA22D0 U7537 ( .A1(n7566), .A2(prog_data[2]), .B1(\mem[252][2] ), .B2(n7565), 
        .Z(n623) );
  OA22D0 U7538 ( .A1(n7566), .A2(prog_data[1]), .B1(\mem[252][1] ), .B2(n7565), 
        .Z(n622) );
  OA22D0 U7539 ( .A1(n7566), .A2(prog_data[0]), .B1(\mem[252][0] ), .B2(n7565), 
        .Z(n621) );
  NR2D0 U7540 ( .A1(n7567), .A2(n7573), .ZN(n7568) );
  INVD0 U7541 ( .I(n7568), .ZN(n7569) );
  OA22D0 U7542 ( .A1(n7569), .A2(prog_data[15]), .B1(\mem[253][15] ), .B2(
        n7568), .Z(n620) );
  OA22D0 U7543 ( .A1(n7569), .A2(prog_data[14]), .B1(\mem[253][14] ), .B2(
        n7568), .Z(n619) );
  OA22D0 U7544 ( .A1(n7569), .A2(prog_data[13]), .B1(\mem[253][13] ), .B2(
        n7568), .Z(n618) );
  OA22D0 U7545 ( .A1(n7569), .A2(prog_data[12]), .B1(\mem[253][12] ), .B2(
        n7568), .Z(n617) );
  OA22D0 U7546 ( .A1(n7569), .A2(prog_data[11]), .B1(\mem[253][11] ), .B2(
        n7568), .Z(n616) );
  OA22D0 U7547 ( .A1(n7569), .A2(prog_data[10]), .B1(\mem[253][10] ), .B2(
        n7568), .Z(n615) );
  OA22D0 U7548 ( .A1(n7569), .A2(prog_data[9]), .B1(\mem[253][9] ), .B2(n7568), 
        .Z(n614) );
  OA22D0 U7549 ( .A1(n7569), .A2(prog_data[8]), .B1(\mem[253][8] ), .B2(n7568), 
        .Z(n613) );
  OA22D0 U7550 ( .A1(n7569), .A2(prog_data[7]), .B1(\mem[253][7] ), .B2(n7568), 
        .Z(n612) );
  OA22D0 U7551 ( .A1(n7569), .A2(prog_data[6]), .B1(\mem[253][6] ), .B2(n7568), 
        .Z(n611) );
  OA22D0 U7552 ( .A1(n7569), .A2(prog_data[5]), .B1(\mem[253][5] ), .B2(n7568), 
        .Z(n610) );
  OA22D0 U7553 ( .A1(n7569), .A2(prog_data[4]), .B1(\mem[253][4] ), .B2(n7568), 
        .Z(n609) );
  OA22D0 U7554 ( .A1(n7569), .A2(prog_data[3]), .B1(\mem[253][3] ), .B2(n7568), 
        .Z(n608) );
  OA22D0 U7555 ( .A1(n7569), .A2(prog_data[2]), .B1(\mem[253][2] ), .B2(n7568), 
        .Z(n607) );
  OA22D0 U7556 ( .A1(n7569), .A2(prog_data[1]), .B1(\mem[253][1] ), .B2(n7568), 
        .Z(n606) );
  OA22D0 U7557 ( .A1(n7569), .A2(prog_data[0]), .B1(\mem[253][0] ), .B2(n7568), 
        .Z(n605) );
  NR2D0 U7558 ( .A1(n7570), .A2(n7573), .ZN(n7571) );
  INVD0 U7559 ( .I(n7571), .ZN(n7572) );
  OA22D0 U7560 ( .A1(n7572), .A2(prog_data[15]), .B1(\mem[254][15] ), .B2(
        n7571), .Z(n604) );
  OA22D0 U7561 ( .A1(n7572), .A2(prog_data[14]), .B1(\mem[254][14] ), .B2(
        n7571), .Z(n603) );
  OA22D0 U7562 ( .A1(n7572), .A2(prog_data[13]), .B1(\mem[254][13] ), .B2(
        n7571), .Z(n602) );
  OA22D0 U7563 ( .A1(n7572), .A2(prog_data[12]), .B1(\mem[254][12] ), .B2(
        n7571), .Z(n601) );
  OA22D0 U7564 ( .A1(n7572), .A2(prog_data[11]), .B1(\mem[254][11] ), .B2(
        n7571), .Z(n600) );
  OA22D0 U7565 ( .A1(n7572), .A2(prog_data[10]), .B1(\mem[254][10] ), .B2(
        n7571), .Z(n599) );
  OA22D0 U7566 ( .A1(n7572), .A2(prog_data[9]), .B1(\mem[254][9] ), .B2(n7571), 
        .Z(n598) );
  OA22D0 U7567 ( .A1(n7572), .A2(prog_data[8]), .B1(\mem[254][8] ), .B2(n7571), 
        .Z(n597) );
  OA22D0 U7568 ( .A1(n7572), .A2(prog_data[7]), .B1(\mem[254][7] ), .B2(n7571), 
        .Z(n596) );
  OA22D0 U7569 ( .A1(n7572), .A2(prog_data[6]), .B1(\mem[254][6] ), .B2(n7571), 
        .Z(n595) );
  OA22D0 U7570 ( .A1(n7572), .A2(prog_data[5]), .B1(\mem[254][5] ), .B2(n7571), 
        .Z(n594) );
  OA22D0 U7571 ( .A1(n7572), .A2(prog_data[4]), .B1(\mem[254][4] ), .B2(n7571), 
        .Z(n593) );
  OA22D0 U7572 ( .A1(n7572), .A2(prog_data[3]), .B1(\mem[254][3] ), .B2(n7571), 
        .Z(n592) );
  OA22D0 U7573 ( .A1(n7572), .A2(prog_data[2]), .B1(\mem[254][2] ), .B2(n7571), 
        .Z(n591) );
  OA22D0 U7574 ( .A1(n7572), .A2(prog_data[1]), .B1(\mem[254][1] ), .B2(n7571), 
        .Z(n590) );
  OA22D0 U7575 ( .A1(n7572), .A2(prog_data[0]), .B1(\mem[254][0] ), .B2(n7571), 
        .Z(n589) );
  NR2D0 U7576 ( .A1(n7574), .A2(n7573), .ZN(n7575) );
  INVD0 U7577 ( .I(n7575), .ZN(n7576) );
  OA22D0 U7578 ( .A1(n7576), .A2(prog_data[15]), .B1(\mem[255][15] ), .B2(
        n7575), .Z(n588) );
  OA22D0 U7579 ( .A1(n7576), .A2(prog_data[14]), .B1(\mem[255][14] ), .B2(
        n7575), .Z(n587) );
  OA22D0 U7580 ( .A1(n7576), .A2(prog_data[13]), .B1(\mem[255][13] ), .B2(
        n7575), .Z(n586) );
  OA22D0 U7581 ( .A1(n7576), .A2(prog_data[12]), .B1(\mem[255][12] ), .B2(
        n7575), .Z(n585) );
  OA22D0 U7582 ( .A1(n7576), .A2(prog_data[11]), .B1(\mem[255][11] ), .B2(
        n7575), .Z(n584) );
  OA22D0 U7583 ( .A1(n7576), .A2(prog_data[10]), .B1(\mem[255][10] ), .B2(
        n7575), .Z(n583) );
  OA22D0 U7584 ( .A1(n7576), .A2(prog_data[9]), .B1(\mem[255][9] ), .B2(n7575), 
        .Z(n582) );
  OA22D0 U7585 ( .A1(n7576), .A2(prog_data[8]), .B1(\mem[255][8] ), .B2(n7575), 
        .Z(n581) );
  OA22D0 U7586 ( .A1(n7576), .A2(prog_data[7]), .B1(\mem[255][7] ), .B2(n7575), 
        .Z(n580) );
  OA22D0 U7587 ( .A1(n7576), .A2(prog_data[6]), .B1(\mem[255][6] ), .B2(n7575), 
        .Z(n579) );
  OA22D0 U7588 ( .A1(n7576), .A2(prog_data[5]), .B1(\mem[255][5] ), .B2(n7575), 
        .Z(n578) );
  OA22D0 U7589 ( .A1(n7576), .A2(prog_data[4]), .B1(\mem[255][4] ), .B2(n7575), 
        .Z(n577) );
  OA22D0 U7590 ( .A1(n7576), .A2(prog_data[3]), .B1(\mem[255][3] ), .B2(n7575), 
        .Z(n576) );
  OA22D0 U7591 ( .A1(n7576), .A2(prog_data[2]), .B1(\mem[255][2] ), .B2(n7575), 
        .Z(n575) );
  OA22D0 U7592 ( .A1(n7576), .A2(prog_data[1]), .B1(\mem[255][1] ), .B2(n7575), 
        .Z(n574) );
  OA22D0 U7593 ( .A1(n7576), .A2(prog_data[0]), .B1(\mem[255][0] ), .B2(n7575), 
        .Z(n573) );
endmodule
