// Created by ihdl
module au ( clk, rst_n, start, R, S, I, ctl_d, result_comb, result_comb_valid, 
        result, done, busy );
  input [23:0] R;
  input [23:0] S;
  input [23:0] I;
  input [1:0] ctl_d;
  output [23:0] result_comb;
  output [23:0] result;
  input clk, rst_n, start;
  output result_comb_valid, done, busy;
  wire   N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, \add_sm[23] , N126, N127,
         N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138,
         N139, N140, N141, N142, N143, N144, N145, N146, N147, N148,
         \sub_sm[23] , \S_lat[23] , \S_mag_safe[0] , inv_start_d, inv_rdy,
         \R_lat[23] , \div_sm[23] , inv_start, N200, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n96, \mult_x_13/n686 , \mult_x_13/n679 ,
         \mult_x_13/n678 , \mult_x_13/n677 , \mult_x_13/n676 ,
         \mult_x_13/n675 , \mult_x_13/n674 , \mult_x_13/n673 ,
         \mult_x_13/n672 , \mult_x_13/n671 , \mult_x_13/n670 ,
         \mult_x_13/n669 , \mult_x_13/n668 , \mult_x_13/n667 ,
         \mult_x_13/n666 , \mult_x_13/n665 , \mult_x_13/n664 ,
         \mult_x_13/n663 , \mult_x_13/n662 , \mult_x_13/n661 ,
         \mult_x_13/n660 , \mult_x_13/n656 , \mult_x_13/n655 ,
         \mult_x_13/n654 , \mult_x_13/n653 , \mult_x_13/n652 ,
         \mult_x_13/n651 , \mult_x_13/n650 , \mult_x_13/n649 ,
         \mult_x_13/n648 , \mult_x_13/n647 , \mult_x_13/n646 ,
         \mult_x_13/n645 , \mult_x_13/n644 , \mult_x_13/n643 ,
         \mult_x_13/n642 , \mult_x_13/n641 , \mult_x_13/n640 ,
         \mult_x_13/n639 , \mult_x_13/n638 , \mult_x_13/n637 ,
         \mult_x_13/n636 , \mult_x_13/n635 , \mult_x_13/n627 ,
         \mult_x_13/n626 , \mult_x_13/n625 , \mult_x_13/n624 ,
         \mult_x_13/n623 , \mult_x_13/n622 , \mult_x_13/n621 ,
         \mult_x_13/n620 , \mult_x_13/n619 , \mult_x_13/n618 ,
         \mult_x_13/n617 , \mult_x_13/n616 , \mult_x_13/n615 ,
         \mult_x_13/n614 , \mult_x_13/n613 , \mult_x_13/n612 ,
         \mult_x_13/n611 , \mult_x_13/n610 , \mult_x_13/n609 ,
         \mult_x_13/n608 , \mult_x_13/n604 , \mult_x_13/n603 ,
         \mult_x_13/n602 , \mult_x_13/n601 , \mult_x_13/n600 ,
         \mult_x_13/n599 , \mult_x_13/n598 , \mult_x_13/n597 ,
         \mult_x_13/n596 , \mult_x_13/n595 , \mult_x_13/n594 ,
         \mult_x_13/n593 , \mult_x_13/n592 , \mult_x_13/n591 ,
         \mult_x_13/n590 , \mult_x_13/n589 , \mult_x_13/n588 ,
         \mult_x_13/n587 , \mult_x_13/n586 , \mult_x_13/n585 ,
         \mult_x_13/n584 , \mult_x_13/n583 , \mult_x_13/n575 ,
         \mult_x_13/n574 , \mult_x_13/n573 , \mult_x_13/n572 ,
         \mult_x_13/n571 , \mult_x_13/n570 , \mult_x_13/n569 ,
         \mult_x_13/n568 , \mult_x_13/n567 , \mult_x_13/n566 ,
         \mult_x_13/n565 , \mult_x_13/n564 , \mult_x_13/n563 ,
         \mult_x_13/n562 , \mult_x_13/n561 , \mult_x_13/n560 ,
         \mult_x_13/n559 , \mult_x_13/n558 , \mult_x_13/n557 ,
         \mult_x_13/n556 , \mult_x_13/n552 , \mult_x_13/n551 ,
         \mult_x_13/n550 , \mult_x_13/n549 , \mult_x_13/n548 ,
         \mult_x_13/n547 , \mult_x_13/n546 , \mult_x_13/n545 ,
         \mult_x_13/n542 , \mult_x_13/n541 , \mult_x_13/n540 ,
         \mult_x_13/n539 , \mult_x_13/n537 , \mult_x_13/n536 ,
         \mult_x_13/n535 , \mult_x_13/n534 , \mult_x_13/n533 ,
         \mult_x_13/n529 , \mult_x_13/n528 , \mult_x_13/n527 ,
         \mult_x_13/n526 , \mult_x_13/n525 , \mult_x_13/n524 ,
         \mult_x_13/n523 , \mult_x_13/n522 , \mult_x_13/n518 ,
         \mult_x_13/n517 , \mult_x_13/n513 , \mult_x_13/n512 ,
         \mult_x_13/n511 , \mult_x_13/n421 , \mult_x_13/n419 ,
         \mult_x_13/n418 , \mult_x_13/n416 , \mult_x_13/n415 ,
         \mult_x_13/n414 , \mult_x_13/n413 , \mult_x_13/n411 ,
         \mult_x_13/n410 , \mult_x_13/n409 , \mult_x_13/n408 ,
         \mult_x_13/n406 , \mult_x_13/n405 , \mult_x_13/n404 ,
         \mult_x_13/n401 , \mult_x_13/n399 , \mult_x_13/n398 ,
         \mult_x_13/n397 , \mult_x_13/n394 , \mult_x_13/n392 ,
         \mult_x_13/n391 , \mult_x_13/n390 , \mult_x_13/n388 ,
         \mult_x_13/n387 , \mult_x_13/n386 , \mult_x_13/n385 ,
         \mult_x_13/n384 , \mult_x_13/n383 , \mult_x_13/n382 ,
         \mult_x_13/n380 , \mult_x_13/n379 , \mult_x_13/n378 ,
         \mult_x_13/n377 , \mult_x_13/n376 , \mult_x_13/n375 ,
         \mult_x_13/n374 , \mult_x_13/n372 , \mult_x_13/n371 ,
         \mult_x_13/n370 , \mult_x_13/n369 , \mult_x_13/n368 ,
         \mult_x_13/n367 , \mult_x_13/n366 , \mult_x_13/n364 ,
         \mult_x_13/n363 , \mult_x_13/n362 , \mult_x_13/n361 ,
         \mult_x_13/n360 , \mult_x_13/n359 , \mult_x_13/n356 ,
         \mult_x_13/n354 , \mult_x_13/n353 , \mult_x_13/n352 ,
         \mult_x_13/n351 , \mult_x_13/n350 , \mult_x_13/n349 ,
         \mult_x_13/n346 , \mult_x_13/n344 , \mult_x_13/n343 ,
         \mult_x_13/n342 , \mult_x_13/n341 , \mult_x_13/n340 ,
         \mult_x_13/n339 , \mult_x_13/n337 , \mult_x_13/n336 ,
         \mult_x_13/n335 , \mult_x_13/n334 , \mult_x_13/n333 ,
         \mult_x_13/n332 , \mult_x_13/n331 , \mult_x_13/n330 ,
         \mult_x_13/n329 , \mult_x_13/n328 , \mult_x_13/n327 ,
         \mult_x_13/n326 , \mult_x_13/n325 , \mult_x_13/n324 ,
         \mult_x_13/n323 , \mult_x_13/n322 , \mult_x_13/n321 ,
         \mult_x_13/n320 , \mult_x_13/n319 , \mult_x_13/n318 ,
         \mult_x_13/n317 , \mult_x_13/n316 , \mult_x_13/n315 ,
         \mult_x_13/n314 , \mult_x_13/n313 , \mult_x_13/n312 ,
         \mult_x_13/n311 , \mult_x_13/n310 , \mult_x_13/n309 ,
         \mult_x_13/n308 , \mult_x_13/n307 , \mult_x_13/n306 ,
         \mult_x_13/n305 , \mult_x_13/n304 , \mult_x_13/n303 ,
         \mult_x_13/n302 , \mult_x_13/n301 , \mult_x_13/n300 ,
         \mult_x_13/n299 , \mult_x_13/n298 , \mult_x_13/n297 ,
         \mult_x_13/n296 , \mult_x_13/n295 , \mult_x_13/n294 ,
         \mult_x_13/n293 , \mult_x_13/n292 , \mult_x_13/n291 ,
         \mult_x_13/n290 , \mult_x_13/n289 , \mult_x_13/n288 ,
         \mult_x_13/n287 , \mult_x_13/n286 , \mult_x_13/n285 ,
         \mult_x_13/n284 , \mult_x_13/n283 , \mult_x_13/n282 ,
         \mult_x_13/n281 , \mult_x_13/n280 , \mult_x_13/n279 ,
         \mult_x_13/n278 , \mult_x_13/n277 , \mult_x_13/n276 ,
         \mult_x_13/n275 , \mult_x_13/n274 , \mult_x_13/n273 ,
         \mult_x_13/n272 , \mult_x_13/n271 , \mult_x_13/n270 ,
         \mult_x_13/n269 , \mult_x_13/n268 , \mult_x_13/n267 ,
         \mult_x_13/n266 , \mult_x_13/n265 , \mult_x_13/n264 ,
         \mult_x_13/n263 , \mult_x_13/n262 , \mult_x_13/n261 ,
         \mult_x_13/n260 , \mult_x_13/n259 , \mult_x_13/n258 ,
         \mult_x_13/n256 , \mult_x_13/n255 , \mult_x_13/n254 ,
         \mult_x_13/n253 , \mult_x_13/n252 , \mult_x_13/n251 ,
         \mult_x_13/n250 , \mult_x_13/n249 , \mult_x_13/n247 ,
         \mult_x_13/n246 , \mult_x_13/n245 , \mult_x_13/n244 ,
         \mult_x_13/n243 , \mult_x_13/n242 , \mult_x_13/n241 ,
         \mult_x_13/n240 , \mult_x_13/n239 , \mult_x_13/n238 ,
         \mult_x_13/n237 , \mult_x_13/n236 , \mult_x_13/n235 ,
         \mult_x_13/n234 , \mult_x_13/n233 , \mult_x_13/n232 ,
         \mult_x_13/n231 , \mult_x_13/n230 , \mult_x_13/n229 ,
         \mult_x_13/n228 , \mult_x_13/n227 , \mult_x_13/n226 ,
         \mult_x_13/n225 , \mult_x_13/n224 , \mult_x_13/n222 ,
         \mult_x_13/n221 , \mult_x_13/n220 , \mult_x_13/n219 ,
         \mult_x_13/n218 , \mult_x_13/n217 , \mult_x_13/n216 ,
         \mult_x_13/n215 , \mult_x_13/n214 , \mult_x_13/n213 ,
         \mult_x_13/n212 , \mult_x_13/n211 , \mult_x_13/n209 ,
         \mult_x_13/n207 , \mult_x_13/n206 , \mult_x_13/n205 ,
         \mult_x_13/n203 , \mult_x_13/n202 , \mult_x_13/n201 ,
         \mult_x_13/n200 , \mult_x_13/n199 , \mult_x_13/n198 ,
         \mult_x_13/n197 , \mult_x_13/n196 , \mult_x_13/n195 ,
         \mult_x_13/n194 , \mult_x_13/n193 , \mult_x_13/n192 ,
         \mult_x_13/n191 , \mult_x_13/n190 , \mult_x_13/n188 ,
         \mult_x_13/n187 , \mult_x_13/n186 , \mult_x_13/n185 ,
         \mult_x_13/n184 , \mult_x_13/n183 , \mult_x_13/n178 , \mult_x_9/n686 ,
         \mult_x_9/n679 , \mult_x_9/n678 , \mult_x_9/n677 , \mult_x_9/n676 ,
         \mult_x_9/n675 , \mult_x_9/n674 , \mult_x_9/n673 , \mult_x_9/n672 ,
         \mult_x_9/n671 , \mult_x_9/n670 , \mult_x_9/n669 , \mult_x_9/n668 ,
         \mult_x_9/n667 , \mult_x_9/n666 , \mult_x_9/n665 , \mult_x_9/n664 ,
         \mult_x_9/n663 , \mult_x_9/n662 , \mult_x_9/n661 , \mult_x_9/n660 ,
         \mult_x_9/n656 , \mult_x_9/n655 , \mult_x_9/n654 , \mult_x_9/n653 ,
         \mult_x_9/n652 , \mult_x_9/n651 , \mult_x_9/n650 , \mult_x_9/n649 ,
         \mult_x_9/n648 , \mult_x_9/n647 , \mult_x_9/n646 , \mult_x_9/n645 ,
         \mult_x_9/n644 , \mult_x_9/n643 , \mult_x_9/n642 , \mult_x_9/n641 ,
         \mult_x_9/n640 , \mult_x_9/n639 , \mult_x_9/n638 , \mult_x_9/n637 ,
         \mult_x_9/n636 , \mult_x_9/n635 , \mult_x_9/n627 , \mult_x_9/n626 ,
         \mult_x_9/n625 , \mult_x_9/n624 , \mult_x_9/n623 , \mult_x_9/n622 ,
         \mult_x_9/n621 , \mult_x_9/n620 , \mult_x_9/n619 , \mult_x_9/n618 ,
         \mult_x_9/n617 , \mult_x_9/n616 , \mult_x_9/n615 , \mult_x_9/n614 ,
         \mult_x_9/n613 , \mult_x_9/n612 , \mult_x_9/n611 , \mult_x_9/n610 ,
         \mult_x_9/n609 , \mult_x_9/n608 , \mult_x_9/n604 , \mult_x_9/n603 ,
         \mult_x_9/n602 , \mult_x_9/n601 , \mult_x_9/n600 , \mult_x_9/n599 ,
         \mult_x_9/n598 , \mult_x_9/n597 , \mult_x_9/n596 , \mult_x_9/n595 ,
         \mult_x_9/n594 , \mult_x_9/n593 , \mult_x_9/n592 , \mult_x_9/n591 ,
         \mult_x_9/n590 , \mult_x_9/n589 , \mult_x_9/n588 , \mult_x_9/n587 ,
         \mult_x_9/n586 , \mult_x_9/n585 , \mult_x_9/n584 , \mult_x_9/n583 ,
         \mult_x_9/n575 , \mult_x_9/n574 , \mult_x_9/n573 , \mult_x_9/n572 ,
         \mult_x_9/n571 , \mult_x_9/n570 , \mult_x_9/n569 , \mult_x_9/n568 ,
         \mult_x_9/n567 , \mult_x_9/n566 , \mult_x_9/n565 , \mult_x_9/n564 ,
         \mult_x_9/n563 , \mult_x_9/n562 , \mult_x_9/n561 , \mult_x_9/n560 ,
         \mult_x_9/n559 , \mult_x_9/n558 , \mult_x_9/n557 , \mult_x_9/n556 ,
         \mult_x_9/n552 , \mult_x_9/n551 , \mult_x_9/n550 , \mult_x_9/n549 ,
         \mult_x_9/n548 , \mult_x_9/n547 , \mult_x_9/n546 , \mult_x_9/n545 ,
         \mult_x_9/n542 , \mult_x_9/n541 , \mult_x_9/n540 , \mult_x_9/n539 ,
         \mult_x_9/n537 , \mult_x_9/n536 , \mult_x_9/n535 , \mult_x_9/n534 ,
         \mult_x_9/n533 , \mult_x_9/n529 , \mult_x_9/n528 , \mult_x_9/n527 ,
         \mult_x_9/n526 , \mult_x_9/n525 , \mult_x_9/n524 , \mult_x_9/n523 ,
         \mult_x_9/n522 , \mult_x_9/n518 , \mult_x_9/n517 , \mult_x_9/n513 ,
         \mult_x_9/n512 , \mult_x_9/n511 , \mult_x_9/n421 , \mult_x_9/n419 ,
         \mult_x_9/n418 , \mult_x_9/n416 , \mult_x_9/n415 , \mult_x_9/n414 ,
         \mult_x_9/n413 , \mult_x_9/n411 , \mult_x_9/n410 , \mult_x_9/n409 ,
         \mult_x_9/n408 , \mult_x_9/n406 , \mult_x_9/n405 , \mult_x_9/n404 ,
         \mult_x_9/n401 , \mult_x_9/n399 , \mult_x_9/n398 , \mult_x_9/n397 ,
         \mult_x_9/n394 , \mult_x_9/n392 , \mult_x_9/n391 , \mult_x_9/n390 ,
         \mult_x_9/n388 , \mult_x_9/n387 , \mult_x_9/n386 , \mult_x_9/n385 ,
         \mult_x_9/n384 , \mult_x_9/n383 , \mult_x_9/n382 , \mult_x_9/n380 ,
         \mult_x_9/n379 , \mult_x_9/n378 , \mult_x_9/n377 , \mult_x_9/n376 ,
         \mult_x_9/n375 , \mult_x_9/n374 , \mult_x_9/n372 , \mult_x_9/n371 ,
         \mult_x_9/n370 , \mult_x_9/n369 , \mult_x_9/n368 , \mult_x_9/n367 ,
         \mult_x_9/n366 , \mult_x_9/n364 , \mult_x_9/n363 , \mult_x_9/n362 ,
         \mult_x_9/n361 , \mult_x_9/n360 , \mult_x_9/n359 , \mult_x_9/n356 ,
         \mult_x_9/n354 , \mult_x_9/n353 , \mult_x_9/n352 , \mult_x_9/n351 ,
         \mult_x_9/n350 , \mult_x_9/n349 , \mult_x_9/n346 , \mult_x_9/n344 ,
         \mult_x_9/n343 , \mult_x_9/n342 , \mult_x_9/n341 , \mult_x_9/n340 ,
         \mult_x_9/n339 , \mult_x_9/n337 , \mult_x_9/n336 , \mult_x_9/n335 ,
         \mult_x_9/n334 , \mult_x_9/n333 , \mult_x_9/n332 , \mult_x_9/n331 ,
         \mult_x_9/n330 , \mult_x_9/n329 , \mult_x_9/n328 , \mult_x_9/n327 ,
         \mult_x_9/n326 , \mult_x_9/n325 , \mult_x_9/n324 , \mult_x_9/n323 ,
         \mult_x_9/n322 , \mult_x_9/n321 , \mult_x_9/n320 , \mult_x_9/n319 ,
         \mult_x_9/n318 , \mult_x_9/n317 , \mult_x_9/n316 , \mult_x_9/n315 ,
         \mult_x_9/n314 , \mult_x_9/n313 , \mult_x_9/n312 , \mult_x_9/n311 ,
         \mult_x_9/n310 , \mult_x_9/n309 , \mult_x_9/n308 , \mult_x_9/n307 ,
         \mult_x_9/n306 , \mult_x_9/n305 , \mult_x_9/n304 , \mult_x_9/n303 ,
         \mult_x_9/n302 , \mult_x_9/n301 , \mult_x_9/n300 , \mult_x_9/n299 ,
         \mult_x_9/n298 , \mult_x_9/n297 , \mult_x_9/n296 , \mult_x_9/n295 ,
         \mult_x_9/n294 , \mult_x_9/n293 , \mult_x_9/n292 , \mult_x_9/n291 ,
         \mult_x_9/n290 , \mult_x_9/n289 , \mult_x_9/n288 , \mult_x_9/n287 ,
         \mult_x_9/n286 , \mult_x_9/n285 , \mult_x_9/n284 , \mult_x_9/n283 ,
         \mult_x_9/n282 , \mult_x_9/n281 , \mult_x_9/n280 , \mult_x_9/n279 ,
         \mult_x_9/n278 , \mult_x_9/n277 , \mult_x_9/n276 , \mult_x_9/n275 ,
         \mult_x_9/n274 , \mult_x_9/n273 , \mult_x_9/n272 , \mult_x_9/n271 ,
         \mult_x_9/n270 , \mult_x_9/n269 , \mult_x_9/n268 , \mult_x_9/n267 ,
         \mult_x_9/n266 , \mult_x_9/n265 , \mult_x_9/n264 , \mult_x_9/n263 ,
         \mult_x_9/n262 , \mult_x_9/n261 , \mult_x_9/n260 , \mult_x_9/n259 ,
         \mult_x_9/n258 , \mult_x_9/n256 , \mult_x_9/n255 , \mult_x_9/n254 ,
         \mult_x_9/n253 , \mult_x_9/n252 , \mult_x_9/n251 , \mult_x_9/n250 ,
         \mult_x_9/n249 , \mult_x_9/n247 , \mult_x_9/n246 , \mult_x_9/n245 ,
         \mult_x_9/n244 , \mult_x_9/n243 , \mult_x_9/n242 , \mult_x_9/n241 ,
         \mult_x_9/n240 , \mult_x_9/n239 , \mult_x_9/n238 , \mult_x_9/n237 ,
         \mult_x_9/n236 , \mult_x_9/n235 , \mult_x_9/n234 , \mult_x_9/n233 ,
         \mult_x_9/n232 , \mult_x_9/n231 , \mult_x_9/n230 , \mult_x_9/n229 ,
         \mult_x_9/n228 , \mult_x_9/n227 , \mult_x_9/n226 , \mult_x_9/n225 ,
         \mult_x_9/n224 , \mult_x_9/n222 , \mult_x_9/n221 , \mult_x_9/n220 ,
         \mult_x_9/n219 , \mult_x_9/n218 , \mult_x_9/n217 , \mult_x_9/n216 ,
         \mult_x_9/n215 , \mult_x_9/n214 , \mult_x_9/n213 , \mult_x_9/n212 ,
         \mult_x_9/n211 , \mult_x_9/n209 , \mult_x_9/n207 , \mult_x_9/n206 ,
         \mult_x_9/n205 , \mult_x_9/n203 , \mult_x_9/n202 , \mult_x_9/n201 ,
         \mult_x_9/n200 , \mult_x_9/n199 , \mult_x_9/n198 , \mult_x_9/n197 ,
         \mult_x_9/n196 , \mult_x_9/n195 , \mult_x_9/n194 , \mult_x_9/n193 ,
         \mult_x_9/n192 , \mult_x_9/n191 , \mult_x_9/n190 , \mult_x_9/n188 ,
         \mult_x_9/n187 , \mult_x_9/n186 , \mult_x_9/n185 , \mult_x_9/n184 ,
         \mult_x_9/n183 , \mult_x_9/n178 , n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267;
  wire   [24:0] add_tc;
  wire   [24:0] sub_tc;
  wire   [45:14] prod_full;
  wire   [22:0] S_lat_mag;
  wire   [22:0] inv_Q_mag;
  wire   [22:0] R_lat_mag;
  wire   [22:0] div_mag_sat;
  wire   [1:0] state;
  wire   [1:0] next_state;

  mult_inv Mult_Inv ( .clk(clk), .rst_n(rst_n), .start(inv_start_d), .S_mag({
        S_lat_mag[22:1], \S_mag_safe[0] }), .Q_mag(inv_Q_mag), .rdy(inv_rdy)
         );
  DFCNQD1 \state_reg[0]  ( .D(next_state[0]), .CP(clk), .CDN(rst_n), .Q(
        state[0]) );
  DFCNQD1 done_reg ( .D(n96), .CP(clk), .CDN(rst_n), .Q(done) );
  DFCNQD1 inv_start_d_reg ( .D(inv_start), .CP(clk), .CDN(rst_n), .Q(
        inv_start_d) );
  DFCNQD1 \state_reg[1]  ( .D(next_state[1]), .CP(clk), .CDN(rst_n), .Q(
        state[1]) );
  EDFQD1 \R_lat_reg[0]  ( .D(R[0]), .E(n2267), .CP(clk), .Q(R_lat_mag[0]) );
  EDFQD1 \S_lat_reg[23]  ( .D(S[23]), .E(n2267), .CP(clk), .Q(\S_lat[23] ) );
  EDFQD1 \S_lat_reg[22]  ( .D(S[22]), .E(n2267), .CP(clk), .Q(S_lat_mag[22])
         );
  EDFQD1 \S_lat_reg[21]  ( .D(S[21]), .E(n2267), .CP(clk), .Q(S_lat_mag[21])
         );
  EDFQD1 \S_lat_reg[20]  ( .D(S[20]), .E(n2267), .CP(clk), .Q(S_lat_mag[20])
         );
  EDFQD1 \S_lat_reg[19]  ( .D(S[19]), .E(n2267), .CP(clk), .Q(S_lat_mag[19])
         );
  EDFQD1 \S_lat_reg[18]  ( .D(S[18]), .E(n2267), .CP(clk), .Q(S_lat_mag[18])
         );
  EDFQD1 \S_lat_reg[17]  ( .D(S[17]), .E(n2267), .CP(clk), .Q(S_lat_mag[17])
         );
  EDFQD1 \S_lat_reg[16]  ( .D(S[16]), .E(n2267), .CP(clk), .Q(S_lat_mag[16])
         );
  EDFQD1 \S_lat_reg[15]  ( .D(S[15]), .E(n2267), .CP(clk), .Q(S_lat_mag[15])
         );
  EDFQD1 \S_lat_reg[14]  ( .D(S[14]), .E(n2267), .CP(clk), .Q(S_lat_mag[14])
         );
  EDFQD1 \S_lat_reg[13]  ( .D(S[13]), .E(n2267), .CP(clk), .Q(S_lat_mag[13])
         );
  EDFQD1 \S_lat_reg[12]  ( .D(S[12]), .E(n2267), .CP(clk), .Q(S_lat_mag[12])
         );
  EDFQD1 \S_lat_reg[11]  ( .D(S[11]), .E(n2267), .CP(clk), .Q(S_lat_mag[11])
         );
  EDFQD1 \S_lat_reg[10]  ( .D(S[10]), .E(n2267), .CP(clk), .Q(S_lat_mag[10])
         );
  EDFQD1 \S_lat_reg[9]  ( .D(S[9]), .E(n2267), .CP(clk), .Q(S_lat_mag[9]) );
  EDFQD1 \S_lat_reg[8]  ( .D(S[8]), .E(n2267), .CP(clk), .Q(S_lat_mag[8]) );
  EDFQD1 \S_lat_reg[7]  ( .D(S[7]), .E(n2267), .CP(clk), .Q(S_lat_mag[7]) );
  EDFQD1 \S_lat_reg[6]  ( .D(S[6]), .E(n2267), .CP(clk), .Q(S_lat_mag[6]) );
  EDFQD1 \S_lat_reg[5]  ( .D(S[5]), .E(n2267), .CP(clk), .Q(S_lat_mag[5]) );
  EDFQD1 \S_lat_reg[4]  ( .D(S[4]), .E(n2267), .CP(clk), .Q(S_lat_mag[4]) );
  EDFQD1 \S_lat_reg[3]  ( .D(S[3]), .E(n2267), .CP(clk), .Q(S_lat_mag[3]) );
  EDFQD1 \S_lat_reg[2]  ( .D(S[2]), .E(n2267), .CP(clk), .Q(S_lat_mag[2]) );
  EDFQD1 \S_lat_reg[1]  ( .D(S[1]), .E(N200), .CP(clk), .Q(S_lat_mag[1]) );
  EDFQD1 \S_lat_reg[0]  ( .D(S[0]), .E(n2267), .CP(clk), .Q(S_lat_mag[0]) );
  EDFQD1 \R_lat_reg[23]  ( .D(R[23]), .E(N200), .CP(clk), .Q(\R_lat[23] ) );
  EDFQD1 \R_lat_reg[22]  ( .D(R[22]), .E(n2267), .CP(clk), .Q(R_lat_mag[22])
         );
  EDFQD1 \R_lat_reg[21]  ( .D(R[21]), .E(N200), .CP(clk), .Q(R_lat_mag[21]) );
  EDFQD1 \R_lat_reg[20]  ( .D(R[20]), .E(n2267), .CP(clk), .Q(R_lat_mag[20])
         );
  EDFQD1 \R_lat_reg[19]  ( .D(R[19]), .E(N200), .CP(clk), .Q(R_lat_mag[19]) );
  EDFQD1 \R_lat_reg[18]  ( .D(R[18]), .E(n2267), .CP(clk), .Q(R_lat_mag[18])
         );
  EDFQD1 \R_lat_reg[17]  ( .D(R[17]), .E(n2267), .CP(clk), .Q(R_lat_mag[17])
         );
  EDFQD1 \R_lat_reg[16]  ( .D(R[16]), .E(n2267), .CP(clk), .Q(R_lat_mag[16])
         );
  EDFQD1 \R_lat_reg[15]  ( .D(R[15]), .E(N200), .CP(clk), .Q(R_lat_mag[15]) );
  EDFQD1 \R_lat_reg[14]  ( .D(R[14]), .E(n2267), .CP(clk), .Q(R_lat_mag[14])
         );
  EDFQD1 \R_lat_reg[13]  ( .D(R[13]), .E(n2267), .CP(clk), .Q(R_lat_mag[13])
         );
  EDFQD1 \R_lat_reg[12]  ( .D(R[12]), .E(n2267), .CP(clk), .Q(R_lat_mag[12])
         );
  EDFQD1 \R_lat_reg[11]  ( .D(R[11]), .E(N200), .CP(clk), .Q(R_lat_mag[11]) );
  EDFQD1 \R_lat_reg[10]  ( .D(R[10]), .E(n2267), .CP(clk), .Q(R_lat_mag[10])
         );
  EDFQD1 \R_lat_reg[9]  ( .D(R[9]), .E(n2267), .CP(clk), .Q(R_lat_mag[9]) );
  EDFQD1 \R_lat_reg[8]  ( .D(R[8]), .E(N200), .CP(clk), .Q(R_lat_mag[8]) );
  EDFQD1 \R_lat_reg[7]  ( .D(R[7]), .E(n2267), .CP(clk), .Q(R_lat_mag[7]) );
  EDFQD1 \R_lat_reg[6]  ( .D(R[6]), .E(N200), .CP(clk), .Q(R_lat_mag[6]) );
  EDFQD1 \R_lat_reg[5]  ( .D(R[5]), .E(N200), .CP(clk), .Q(R_lat_mag[5]) );
  EDFQD1 \R_lat_reg[4]  ( .D(R[4]), .E(n2267), .CP(clk), .Q(R_lat_mag[4]) );
  EDFQD1 \R_lat_reg[3]  ( .D(R[3]), .E(n2267), .CP(clk), .Q(R_lat_mag[3]) );
  EDFQD1 \R_lat_reg[2]  ( .D(R[2]), .E(N200), .CP(clk), .Q(R_lat_mag[2]) );
  EDFQD1 \R_lat_reg[1]  ( .D(R[1]), .E(n2267), .CP(clk), .Q(R_lat_mag[1]) );
  EDFQD1 \result_reg[1]  ( .D(div_mag_sat[1]), .E(n96), .CP(clk), .Q(result[1]) );
  EDFQD1 \result_reg[2]  ( .D(div_mag_sat[2]), .E(n96), .CP(clk), .Q(result[2]) );
  EDFQD1 \result_reg[3]  ( .D(div_mag_sat[3]), .E(n96), .CP(clk), .Q(result[3]) );
  EDFQD1 \result_reg[4]  ( .D(div_mag_sat[4]), .E(n96), .CP(clk), .Q(result[4]) );
  EDFQD1 \result_reg[5]  ( .D(div_mag_sat[5]), .E(n96), .CP(clk), .Q(result[5]) );
  EDFQD1 \result_reg[6]  ( .D(div_mag_sat[6]), .E(n96), .CP(clk), .Q(result[6]) );
  EDFQD1 \result_reg[7]  ( .D(div_mag_sat[7]), .E(n96), .CP(clk), .Q(result[7]) );
  EDFQD1 \result_reg[8]  ( .D(div_mag_sat[8]), .E(n96), .CP(clk), .Q(result[8]) );
  EDFQD1 \result_reg[9]  ( .D(div_mag_sat[9]), .E(n96), .CP(clk), .Q(result[9]) );
  EDFQD1 \result_reg[10]  ( .D(div_mag_sat[10]), .E(n96), .CP(clk), .Q(
        result[10]) );
  EDFQD1 \result_reg[11]  ( .D(div_mag_sat[11]), .E(n96), .CP(clk), .Q(
        result[11]) );
  EDFQD1 \result_reg[12]  ( .D(div_mag_sat[12]), .E(n96), .CP(clk), .Q(
        result[12]) );
  EDFQD1 \result_reg[13]  ( .D(div_mag_sat[13]), .E(n96), .CP(clk), .Q(
        result[13]) );
  EDFQD1 \result_reg[14]  ( .D(div_mag_sat[14]), .E(n96), .CP(clk), .Q(
        result[14]) );
  EDFQD1 \result_reg[15]  ( .D(div_mag_sat[15]), .E(n96), .CP(clk), .Q(
        result[15]) );
  EDFQD1 \result_reg[16]  ( .D(div_mag_sat[16]), .E(n96), .CP(clk), .Q(
        result[16]) );
  EDFQD1 \result_reg[17]  ( .D(div_mag_sat[17]), .E(n96), .CP(clk), .Q(
        result[17]) );
  EDFQD1 \result_reg[18]  ( .D(div_mag_sat[18]), .E(n96), .CP(clk), .Q(
        result[18]) );
  EDFQD1 \result_reg[19]  ( .D(div_mag_sat[19]), .E(n96), .CP(clk), .Q(
        result[19]) );
  EDFQD1 \result_reg[20]  ( .D(div_mag_sat[20]), .E(n96), .CP(clk), .Q(
        result[20]) );
  EDFQD1 \result_reg[21]  ( .D(div_mag_sat[21]), .E(n96), .CP(clk), .Q(
        result[21]) );
  EDFQD1 \result_reg[22]  ( .D(div_mag_sat[22]), .E(n96), .CP(clk), .Q(
        result[22]) );
  EDFQD1 \result_reg[23]  ( .D(\div_sm[23] ), .E(n96), .CP(clk), .Q(result[23]) );
  EDFQD1 \result_reg[0]  ( .D(div_mag_sat[0]), .E(n96), .CP(clk), .Q(result[0]) );
  OR4D0 U5 ( .A1(prod_full[41]), .A2(prod_full[42]), .A3(prod_full[43]), .A4(
        prod_full[44]), .Z(n1) );
  OR4D0 U6 ( .A1(prod_full[39]), .A2(prod_full[37]), .A3(prod_full[45]), .A4(
        n1), .Z(n2) );
  OAI31D0 U8 ( .A1(prod_full[38]), .A2(prod_full[40]), .A3(n2), .B(n79), .ZN(
        n5) );
  OAI221D0 U11 ( .A1(\sub_sm[23] ), .A2(sub_tc[23]), .B1(n69), .B2(N148), .C(
        n78), .ZN(n4) );
  OAI221D0 U14 ( .A1(\add_sm[23] ), .A2(add_tc[23]), .B1(n70), .B2(N97), .C(
        n77), .ZN(n3) );
  CKND2D0 U17 ( .A1(n79), .A2(prod_full[36]), .ZN(n8) );
  OAI221D0 U18 ( .A1(\sub_sm[23] ), .A2(sub_tc[22]), .B1(n69), .B2(N147), .C(
        n78), .ZN(n7) );
  OAI221D0 U19 ( .A1(\add_sm[23] ), .A2(add_tc[22]), .B1(n70), .B2(N96), .C(
        n77), .ZN(n6) );
  ND4D0 U20 ( .A1(n74), .A2(n8), .A3(n7), .A4(n6), .ZN(result_comb[22]) );
  CKND2D0 U21 ( .A1(n79), .A2(prod_full[35]), .ZN(n11) );
  OAI221D0 U22 ( .A1(\sub_sm[23] ), .A2(sub_tc[21]), .B1(n69), .B2(N146), .C(
        n78), .ZN(n10) );
  OAI221D0 U23 ( .A1(\add_sm[23] ), .A2(add_tc[21]), .B1(n70), .B2(N95), .C(
        n77), .ZN(n9) );
  ND4D0 U24 ( .A1(n74), .A2(n11), .A3(n10), .A4(n9), .ZN(result_comb[21]) );
  CKND2D0 U25 ( .A1(n79), .A2(prod_full[34]), .ZN(n14) );
  OAI221D0 U26 ( .A1(\sub_sm[23] ), .A2(sub_tc[20]), .B1(n69), .B2(N145), .C(
        n78), .ZN(n13) );
  OAI221D0 U27 ( .A1(\add_sm[23] ), .A2(add_tc[20]), .B1(n70), .B2(N94), .C(
        n77), .ZN(n12) );
  ND4D0 U28 ( .A1(n74), .A2(n14), .A3(n13), .A4(n12), .ZN(result_comb[20]) );
  CKND2D0 U29 ( .A1(n79), .A2(prod_full[33]), .ZN(n17) );
  OAI221D0 U30 ( .A1(\sub_sm[23] ), .A2(sub_tc[19]), .B1(n69), .B2(N144), .C(
        n78), .ZN(n16) );
  OAI221D0 U31 ( .A1(\add_sm[23] ), .A2(add_tc[19]), .B1(n70), .B2(N93), .C(
        n77), .ZN(n15) );
  CKND2D0 U33 ( .A1(n79), .A2(prod_full[32]), .ZN(n20) );
  OAI221D0 U34 ( .A1(\sub_sm[23] ), .A2(sub_tc[18]), .B1(n69), .B2(N143), .C(
        n78), .ZN(n19) );
  OAI221D0 U35 ( .A1(\add_sm[23] ), .A2(add_tc[18]), .B1(n70), .B2(N92), .C(
        n77), .ZN(n18) );
  ND4D0 U36 ( .A1(n74), .A2(n20), .A3(n19), .A4(n18), .ZN(result_comb[18]) );
  CKND2D0 U37 ( .A1(n79), .A2(prod_full[31]), .ZN(n23) );
  OAI221D0 U38 ( .A1(\sub_sm[23] ), .A2(sub_tc[17]), .B1(n69), .B2(N142), .C(
        n78), .ZN(n22) );
  OAI221D0 U39 ( .A1(\add_sm[23] ), .A2(add_tc[17]), .B1(n70), .B2(N91), .C(
        n77), .ZN(n21) );
  ND4D0 U40 ( .A1(n74), .A2(n23), .A3(n22), .A4(n21), .ZN(result_comb[17]) );
  CKND2D0 U41 ( .A1(n79), .A2(prod_full[30]), .ZN(n26) );
  OAI221D0 U42 ( .A1(\sub_sm[23] ), .A2(sub_tc[16]), .B1(n69), .B2(N141), .C(
        n78), .ZN(n25) );
  OAI221D0 U43 ( .A1(\add_sm[23] ), .A2(add_tc[16]), .B1(n70), .B2(N90), .C(
        n77), .ZN(n24) );
  ND4D0 U44 ( .A1(n74), .A2(n26), .A3(n25), .A4(n24), .ZN(result_comb[16]) );
  CKND2D0 U45 ( .A1(n79), .A2(prod_full[29]), .ZN(n29) );
  OAI221D0 U46 ( .A1(\sub_sm[23] ), .A2(sub_tc[15]), .B1(n69), .B2(N140), .C(
        n78), .ZN(n28) );
  OAI221D0 U47 ( .A1(\add_sm[23] ), .A2(add_tc[15]), .B1(n70), .B2(N89), .C(
        n77), .ZN(n27) );
  CKND2D0 U49 ( .A1(n79), .A2(prod_full[28]), .ZN(n32) );
  OAI221D0 U50 ( .A1(\sub_sm[23] ), .A2(sub_tc[14]), .B1(n69), .B2(N139), .C(
        n78), .ZN(n31) );
  OAI221D0 U51 ( .A1(\add_sm[23] ), .A2(add_tc[14]), .B1(n70), .B2(N88), .C(
        n77), .ZN(n30) );
  ND4D0 U52 ( .A1(n74), .A2(n32), .A3(n31), .A4(n30), .ZN(result_comb[14]) );
  CKND2D0 U53 ( .A1(n79), .A2(prod_full[27]), .ZN(n35) );
  OAI221D0 U54 ( .A1(\sub_sm[23] ), .A2(sub_tc[13]), .B1(n69), .B2(N138), .C(
        n78), .ZN(n34) );
  OAI221D0 U55 ( .A1(\add_sm[23] ), .A2(add_tc[13]), .B1(n70), .B2(N87), .C(
        n77), .ZN(n33) );
  CKND2D0 U57 ( .A1(n79), .A2(prod_full[26]), .ZN(n38) );
  OAI221D0 U58 ( .A1(\sub_sm[23] ), .A2(sub_tc[12]), .B1(n69), .B2(N137), .C(
        n78), .ZN(n37) );
  OAI221D0 U59 ( .A1(\add_sm[23] ), .A2(add_tc[12]), .B1(n70), .B2(N86), .C(
        n77), .ZN(n36) );
  CKND2D0 U61 ( .A1(n79), .A2(prod_full[25]), .ZN(n41) );
  OAI221D0 U62 ( .A1(\sub_sm[23] ), .A2(sub_tc[11]), .B1(n69), .B2(N136), .C(
        n78), .ZN(n40) );
  OAI221D0 U63 ( .A1(\add_sm[23] ), .A2(add_tc[11]), .B1(n70), .B2(N85), .C(
        n77), .ZN(n39) );
  CKND2D0 U65 ( .A1(n79), .A2(prod_full[24]), .ZN(n44) );
  OAI221D0 U66 ( .A1(\sub_sm[23] ), .A2(sub_tc[10]), .B1(n69), .B2(N135), .C(
        n78), .ZN(n43) );
  OAI221D0 U67 ( .A1(\add_sm[23] ), .A2(add_tc[10]), .B1(n70), .B2(N84), .C(
        n77), .ZN(n42) );
  CKND2D0 U69 ( .A1(n79), .A2(prod_full[23]), .ZN(n47) );
  OAI221D0 U70 ( .A1(\sub_sm[23] ), .A2(sub_tc[9]), .B1(n69), .B2(N134), .C(
        n78), .ZN(n46) );
  OAI221D0 U71 ( .A1(\add_sm[23] ), .A2(add_tc[9]), .B1(n70), .B2(N83), .C(n77), .ZN(n45) );
  CKND2D0 U73 ( .A1(n79), .A2(prod_full[22]), .ZN(n50) );
  OAI221D0 U74 ( .A1(\sub_sm[23] ), .A2(sub_tc[8]), .B1(n69), .B2(N133), .C(
        n78), .ZN(n49) );
  OAI221D0 U75 ( .A1(\add_sm[23] ), .A2(add_tc[8]), .B1(n70), .B2(N82), .C(n77), .ZN(n48) );
  CKND2D0 U77 ( .A1(n79), .A2(prod_full[21]), .ZN(n53) );
  OAI221D0 U78 ( .A1(\sub_sm[23] ), .A2(sub_tc[7]), .B1(n69), .B2(N132), .C(
        n78), .ZN(n52) );
  OAI221D0 U79 ( .A1(\add_sm[23] ), .A2(add_tc[7]), .B1(n70), .B2(N81), .C(n77), .ZN(n51) );
  CKND2D0 U81 ( .A1(n79), .A2(prod_full[20]), .ZN(n56) );
  OAI221D0 U82 ( .A1(\sub_sm[23] ), .A2(sub_tc[6]), .B1(n69), .B2(N131), .C(
        n78), .ZN(n55) );
  OAI221D0 U83 ( .A1(\add_sm[23] ), .A2(add_tc[6]), .B1(n70), .B2(N80), .C(n77), .ZN(n54) );
  CKND2D0 U85 ( .A1(n79), .A2(prod_full[19]), .ZN(n59) );
  OAI221D0 U86 ( .A1(\sub_sm[23] ), .A2(sub_tc[5]), .B1(n69), .B2(N130), .C(
        n78), .ZN(n58) );
  OAI221D0 U87 ( .A1(\add_sm[23] ), .A2(add_tc[5]), .B1(n70), .B2(N79), .C(n77), .ZN(n57) );
  CKND2D0 U89 ( .A1(n79), .A2(prod_full[18]), .ZN(n62) );
  OAI221D0 U90 ( .A1(\sub_sm[23] ), .A2(sub_tc[4]), .B1(n69), .B2(N129), .C(
        n78), .ZN(n61) );
  OAI221D0 U91 ( .A1(\add_sm[23] ), .A2(add_tc[4]), .B1(n70), .B2(N78), .C(n77), .ZN(n60) );
  CKND2D0 U93 ( .A1(n79), .A2(prod_full[17]), .ZN(n65) );
  OAI221D0 U94 ( .A1(\sub_sm[23] ), .A2(sub_tc[3]), .B1(n69), .B2(N128), .C(
        n78), .ZN(n64) );
  OAI221D0 U95 ( .A1(\add_sm[23] ), .A2(add_tc[3]), .B1(n70), .B2(N77), .C(n77), .ZN(n63) );
  CKND2D0 U97 ( .A1(n79), .A2(prod_full[16]), .ZN(n68) );
  OAI221D0 U98 ( .A1(\sub_sm[23] ), .A2(sub_tc[2]), .B1(n69), .B2(N127), .C(
        n78), .ZN(n67) );
  OAI221D0 U99 ( .A1(\add_sm[23] ), .A2(add_tc[2]), .B1(n70), .B2(N76), .C(n77), .ZN(n66) );
  CKND2D0 U101 ( .A1(n79), .A2(prod_full[15]), .ZN(n73) );
  OAI221D0 U102 ( .A1(\sub_sm[23] ), .A2(sub_tc[1]), .B1(n69), .B2(N126), .C(
        n78), .ZN(n72) );
  OAI221D0 U103 ( .A1(\add_sm[23] ), .A2(add_tc[1]), .B1(n70), .B2(N75), .C(
        n77), .ZN(n71) );
  AO22D0 U105 ( .A1(n78), .A2(add_tc[0]), .B1(n77), .B2(add_tc[0]), .Z(n75) );
  AO211D0 U106 ( .A1(n79), .A2(prod_full[14]), .B(n76), .C(n75), .Z(
        result_comb[0]) );
  OA222D0 U3 ( .A1(n1728), .A2(n1822), .B1(n1826), .B2(n1418), .C1(n1740), 
        .C2(n1420), .Z(n80) );
  OAI22D0 U4 ( .A1(n1726), .A2(n1151), .B1(n1728), .B2(n1153), .ZN(n1054) );
  OAI22D0 U7 ( .A1(n1825), .A2(n1151), .B1(n1730), .B2(n1153), .ZN(n1063) );
  AOI211D0 U9 ( .A1(n1733), .A2(n1157), .B(n1055), .C(n1054), .ZN(n1057) );
  OAI22D0 U10 ( .A1(n1730), .A2(n1826), .B1(n1726), .B2(n1824), .ZN(n530) );
  NR2D0 U12 ( .A1(n1825), .A2(n1822), .ZN(n531) );
  OAI22D0 U13 ( .A1(n1825), .A2(n1826), .B1(n1730), .B2(n1824), .ZN(n533) );
  OAI22D0 U15 ( .A1(n1817), .A2(n1151), .B1(n1823), .B2(n1153), .ZN(n1088) );
  NR2D0 U16 ( .A1(n1797), .A2(n1470), .ZN(n1009) );
  AOI22D0 U32 ( .A1(n250), .A2(inv_Q_mag[6]), .B1(n251), .B2(inv_Q_mag[7]), 
        .ZN(n151) );
  INVD0 U48 ( .I(n1475), .ZN(n1037) );
  AOI211D0 U56 ( .A1(n1157), .A2(n1815), .B(n1089), .C(n1088), .ZN(n1090) );
  NR2D0 U60 ( .A1(n1823), .A2(n1529), .ZN(n1533) );
  OAI22D0 U64 ( .A1(n1807), .A2(n1531), .B1(n1812), .B2(n1530), .ZN(n1517) );
  NR2D0 U68 ( .A1(n1812), .A2(n1417), .ZN(n1013) );
  AOI22D0 U72 ( .A1(n2256), .A2(inv_Q_mag[4]), .B1(n2255), .B2(n2254), .ZN(
        n2260) );
  OAI22D0 U76 ( .A1(n1757), .A2(n1419), .B1(n1762), .B2(n1394), .ZN(n1035) );
  OAI22D0 U80 ( .A1(n1762), .A2(n1472), .B1(n1767), .B2(n1471), .ZN(n1431) );
  NR2D0 U84 ( .A1(n515), .A2(n516), .ZN(\mult_x_9/n421 ) );
  OAI22D0 U88 ( .A1(n1825), .A2(n1657), .B1(n1730), .B2(n1656), .ZN(n474) );
  NR2D0 U92 ( .A1(n1812), .A2(n1655), .ZN(n1650) );
  NR2D0 U96 ( .A1(n1823), .A2(n1596), .ZN(n1585) );
  CKND2D0 U100 ( .A1(R[20]), .A2(n426), .ZN(n425) );
  AOI211D0 U104 ( .A1(n1475), .A2(n1719), .B(n1465), .C(n1464), .ZN(n1466) );
  NR2D0 U107 ( .A1(n1797), .A2(n1596), .ZN(n1570) );
  OAI22D0 U108 ( .A1(\mult_x_9/n660 ), .A2(R[4]), .B1(n596), .B2(R[5]), .ZN(
        n519) );
  CKND2D0 U109 ( .A1(n1831), .A2(n1385), .ZN(n989) );
  NR2D0 U110 ( .A1(n1787), .A2(n1472), .ZN(n1444) );
  OAI22D0 U111 ( .A1(n1787), .A2(n1419), .B1(n1792), .B2(n1394), .ZN(n941) );
  NR2D0 U112 ( .A1(n1777), .A2(n1417), .ZN(n945) );
  CKND2D0 U113 ( .A1(n1373), .A2(n1372), .ZN(n1374) );
  CKND2D0 U114 ( .A1(n170), .A2(n169), .ZN(n171) );
  AOI211D0 U115 ( .A1(n1385), .A2(n1755), .B(n1036), .C(n1035), .ZN(n1159) );
  OAI22D0 U116 ( .A1(n1747), .A2(n1419), .B1(n1752), .B2(n1394), .ZN(n1026) );
  OAI211D0 U117 ( .A1(n1417), .A2(n1772), .B(n1382), .C(n1381), .ZN(n1410) );
  OAI22D0 U118 ( .A1(n1823), .A2(n1729), .B1(n1825), .B2(n1727), .ZN(n1714) );
  AOI211D0 U119 ( .A1(n1660), .A2(n1719), .B(n475), .C(n474), .ZN(n476) );
  NR2D0 U120 ( .A1(n1807), .A2(n1725), .ZN(n1703) );
  OAI22D0 U121 ( .A1(n1792), .A2(n1729), .B1(n1802), .B2(n1727), .ZN(n1696) );
  NR2D0 U122 ( .A1(n1767), .A2(n1822), .ZN(n1769) );
  NR2D0 U123 ( .A1(n1418), .A2(n1379), .ZN(\mult_x_9/n529 ) );
  AOI211D0 U124 ( .A1(n1785), .A2(n1660), .B(n1632), .C(n1631), .ZN(n1633) );
  OAI211D0 U125 ( .A1(n1417), .A2(n1825), .B(n982), .C(n981), .ZN(
        \mult_x_9/n525 ) );
  OAI22D0 U126 ( .A1(n1772), .A2(n1657), .B1(n1777), .B2(n1656), .ZN(n1622) );
  OAI22D0 U127 ( .A1(n1757), .A2(n1657), .B1(n1762), .B2(n1656), .ZN(n1613) );
  NR2D0 U128 ( .A1(n1767), .A2(n1596), .ZN(n1552) );
  OAI22D0 U129 ( .A1(n1747), .A2(n1598), .B1(n1757), .B2(n1597), .ZN(n1542) );
  AOI22D0 U130 ( .A1(S[11]), .A2(n1384), .B1(S[10]), .B2(n1383), .ZN(n1001) );
  INVD0 U131 ( .I(n1601), .ZN(n1537) );
  AOI211D0 U132 ( .A1(n2178), .A2(n2167), .B(n2166), .C(n2165), .ZN(n2168) );
  AOI22D0 U133 ( .A1(inv_Q_mag[4]), .A2(n1957), .B1(inv_Q_mag[5]), .B2(n1956), 
        .ZN(n503) );
  INVD0 U134 ( .I(\mult_x_9/n183 ), .ZN(n1277) );
  OAI211D0 U135 ( .A1(n1417), .A2(n1762), .B(n963), .C(n962), .ZN(
        \mult_x_9/n512 ) );
  INVD0 U136 ( .I(\mult_x_9/n411 ), .ZN(n1103) );
  OAI22D0 U137 ( .A1(n1817), .A2(n1729), .B1(n1827), .B2(n1727), .ZN(n1711) );
  NR2D0 U138 ( .A1(n1399), .A2(n1317), .ZN(\mult_x_9/n366 ) );
  INVD0 U139 ( .I(n1343), .ZN(\mult_x_9/n336 ) );
  AOI211D0 U140 ( .A1(n1750), .A2(n1830), .B(n1749), .C(n1748), .ZN(n1751) );
  AOI211D0 U141 ( .A1(n1770), .A2(n1660), .B(n1623), .C(n1622), .ZN(n1624) );
  INVD0 U142 ( .I(n1014), .ZN(\mult_x_9/n256 ) );
  INVD0 U143 ( .I(n1313), .ZN(\mult_x_9/n237 ) );
  AOI211D0 U144 ( .A1(n1755), .A2(n1534), .B(n1488), .C(n1487), .ZN(n1489) );
  INVD0 U145 ( .I(\mult_x_13/n416 ), .ZN(n181) );
  AOI22D0 U146 ( .A1(inv_Q_mag[4]), .A2(n2085), .B1(inv_Q_mag[5]), .B2(n2084), 
        .ZN(n564) );
  AOI22D0 U147 ( .A1(inv_Q_mag[7]), .A2(n1955), .B1(n2242), .B2(n1954), .ZN(
        n1946) );
  NR2D0 U148 ( .A1(n2172), .A2(n1893), .ZN(n1897) );
  NR2D0 U149 ( .A1(n2174), .A2(n2021), .ZN(n542) );
  INVD0 U150 ( .I(n1385), .ZN(n1421) );
  INVD0 U151 ( .I(\mult_x_9/n191 ), .ZN(n1280) );
  OAI22D0 U152 ( .A1(n1777), .A2(n1151), .B1(n1782), .B2(n1153), .ZN(n1129) );
  NR2D0 U153 ( .A1(R[0]), .A2(R[1]), .ZN(n1047) );
  NR2D0 U154 ( .A1(S[4]), .A2(n606), .ZN(n592) );
  CKND2D0 U155 ( .A1(n661), .A2(n1736), .ZN(n691) );
  CKAN2D0 U156 ( .A1(n698), .A2(n700), .Z(n707) );
  CKND2D0 U157 ( .A1(n712), .A2(n1787), .ZN(n734) );
  CKAN2D0 U158 ( .A1(n749), .A2(n751), .Z(n761) );
  CKND2D0 U159 ( .A1(n766), .A2(n1477), .ZN(n771) );
  NR2D0 U160 ( .A1(n1408), .A2(n1367), .ZN(\mult_x_13/n408 ) );
  NR2D0 U161 ( .A1(n2127), .A2(n1285), .ZN(n959) );
  AOI22D0 U162 ( .A1(inv_Q_mag[14]), .A2(n1957), .B1(inv_Q_mag[13]), .B2(n1955), .ZN(n1927) );
  AOI22D0 U163 ( .A1(inv_Q_mag[14]), .A2(n2083), .B1(n2214), .B2(n2082), .ZN(
        n2053) );
  AOI22D0 U164 ( .A1(inv_Q_mag[2]), .A2(n1336), .B1(n2177), .B2(n1334), .ZN(
        n1290) );
  CKND2D0 U165 ( .A1(n1952), .A2(n1951), .ZN(n1953) );
  AOI22D0 U166 ( .A1(inv_Q_mag[9]), .A2(n2083), .B1(n2234), .B2(n2082), .ZN(
        n2068) );
  OAI22D0 U167 ( .A1(n2164), .A2(n2023), .B1(n2155), .B2(n2022), .ZN(n2012) );
  AOI22D0 U168 ( .A1(inv_Q_mag[5]), .A2(n2083), .B1(n2250), .B2(n2082), .ZN(
        n2080) );
  INVD0 U169 ( .I(inv_Q_mag[9]), .ZN(n2143) );
  INVD0 U170 ( .I(n1162), .ZN(prod_full[44]) );
  INVD0 U171 ( .I(\mult_x_9/n184 ), .ZN(n1176) );
  INVD0 U172 ( .I(n1359), .ZN(\mult_x_9/n394 ) );
  AOI211D0 U173 ( .A1(n1770), .A2(n1157), .B(n1133), .C(n1132), .ZN(n1134) );
  INVD0 U174 ( .I(S[7]), .ZN(n1817) );
  NR2D0 U175 ( .A1(n714), .A2(n1389), .ZN(n710) );
  CKND2D0 U176 ( .A1(S[23]), .A2(n752), .ZN(n753) );
  NR2D0 U177 ( .A1(n763), .A2(n1389), .ZN(n764) );
  INVD0 U178 ( .I(R[21]), .ZN(n768) );
  NR2D0 U179 ( .A1(n2123), .A2(n1895), .ZN(n1864) );
  AOI22D0 U180 ( .A1(inv_Q_mag[15]), .A2(n1955), .B1(n2210), .B2(n1954), .ZN(
        n1922) );
  OAI22D0 U181 ( .A1(n2103), .A2(n2022), .B1(n2111), .B2(n2023), .ZN(n1973) );
  OAI22D0 U182 ( .A1(n2119), .A2(n2022), .B1(n2123), .B2(n2021), .ZN(n1985) );
  INVD0 U183 ( .I(inv_Q_mag[7]), .ZN(n2151) );
  INVD0 U184 ( .I(n105), .ZN(n99) );
  AOI22D0 U185 ( .A1(inv_Q_mag[20]), .A2(n2256), .B1(n2190), .B2(n2255), .ZN(
        n2192) );
  OAI211D0 U186 ( .A1(n1840), .A2(n2172), .B(n1290), .C(n1289), .ZN(
        \mult_x_13/n526 ) );
  CKND2D0 U187 ( .A1(n2062), .A2(n2061), .ZN(n2063) );
  CKAN2D0 U188 ( .A1(n1380), .A2(inv_Q_mag[0]), .Z(\mult_x_13/n529 ) );
  AOI22D0 U189 ( .A1(inv_Q_mag[14]), .A2(n2257), .B1(inv_Q_mag[13]), .B2(n2256), .ZN(n2219) );
  CKND2D0 U190 ( .A1(n2077), .A2(n2076), .ZN(n2078) );
  INVD0 U191 ( .I(\mult_x_13/n191 ), .ZN(n282) );
  NR2D0 U192 ( .A1(n2107), .A2(n1285), .ZN(n213) );
  NR2D0 U193 ( .A1(n2147), .A2(n2169), .ZN(n2145) );
  INVD0 U194 ( .I(add_tc[23]), .ZN(n2263) );
  INVD0 U195 ( .I(\mult_x_9/n377 ), .ZN(n1213) );
  INVD0 U196 ( .I(\mult_x_9/n351 ), .ZN(n1201) );
  INVD0 U197 ( .I(\mult_x_9/n322 ), .ZN(n1249) );
  AOI32D0 U198 ( .A1(n1157), .A2(\mult_x_9/n686 ), .A3(n1156), .B1(R[2]), .B2(
        n1155), .ZN(n1203) );
  INVD0 U199 ( .I(\mult_x_9/n276 ), .ZN(n1216) );
  INVD0 U200 ( .I(\mult_x_9/n250 ), .ZN(n1268) );
  INVD0 U201 ( .I(\mult_x_9/n225 ), .ZN(n1196) );
  INVD0 U202 ( .I(n798), .ZN(n836) );
  INVD0 U203 ( .I(n1363), .ZN(\mult_x_13/n394 ) );
  OAI22D0 U204 ( .A1(n2185), .A2(n2022), .B1(n2099), .B2(n2023), .ZN(n1964) );
  CKND2D0 U205 ( .A1(n1380), .A2(n211), .ZN(n1840) );
  CKND2D0 U206 ( .A1(n2035), .A2(n2034), .ZN(n2036) );
  CKND2D0 U207 ( .A1(n1931), .A2(n1930), .ZN(n1932) );
  AOI22D0 U208 ( .A1(inv_Q_mag[22]), .A2(n2256), .B1(n2181), .B2(n2255), .ZN(
        n2182) );
  AOI211D0 U209 ( .A1(n2178), .A2(n2202), .B(n2105), .C(n2104), .ZN(n2106) );
  CKND2D0 U210 ( .A1(n2204), .A2(n2203), .ZN(n2205) );
  INVD0 U211 ( .I(n1347), .ZN(\mult_x_13/n336 ) );
  CKND2D0 U212 ( .A1(n2224), .A2(n2223), .ZN(n2225) );
  INVD0 U213 ( .I(n288), .ZN(n298) );
  INVD0 U214 ( .I(n2089), .ZN(n2181) );
  CKND2D0 U215 ( .A1(n262), .A2(n261), .ZN(n274) );
  INVD0 U216 ( .I(R[0]), .ZN(n1046) );
  INVD0 U217 ( .I(n807), .ZN(n642) );
  INVD0 U218 ( .I(n678), .ZN(n679) );
  CKND2D0 U219 ( .A1(n911), .A2(n913), .ZN(n923) );
  NR2D0 U220 ( .A1(sub_tc[8]), .A2(n638), .ZN(n870) );
  INVD0 U221 ( .I(n863), .ZN(n862) );
  INVD0 U222 ( .I(n859), .ZN(n860) );
  INVD0 U223 ( .I(n756), .ZN(n716) );
  INVD0 U224 ( .I(n787), .ZN(n788) );
  NR2D0 U225 ( .A1(sub_tc[18]), .A2(n918), .ZN(n917) );
  INVD0 U226 ( .I(n889), .ZN(n888) );
  INVD0 U227 ( .I(n799), .ZN(n773) );
  CKND2D0 U228 ( .A1(n1913), .A2(n1912), .ZN(n1914) );
  AOI211D0 U229 ( .A1(n2026), .A2(n2198), .B(n1971), .C(n1970), .ZN(n1972) );
  CKND2D0 U230 ( .A1(n2041), .A2(n2040), .ZN(n2042) );
  AOI211D0 U231 ( .A1(n2178), .A2(n2198), .B(n2101), .C(n2100), .ZN(n2102) );
  CKND2D0 U232 ( .A1(inv_Q_mag[22]), .A2(n217), .ZN(n2089) );
  AOI22D0 U233 ( .A1(inv_Q_mag[21]), .A2(n251), .B1(n250), .B2(inv_Q_mag[20]), 
        .ZN(n245) );
  AOI22D0 U234 ( .A1(n250), .A2(inv_Q_mag[18]), .B1(n251), .B2(inv_Q_mag[19]), 
        .ZN(n238) );
  INVD0 U235 ( .I(n280), .ZN(n301) );
  OAI21D0 U236 ( .A1(n262), .A2(n261), .B(n274), .ZN(n272) );
  OAI21D0 U237 ( .A1(S[0]), .A2(n1046), .B(n641), .ZN(add_tc[0]) );
  AOI21D0 U238 ( .A1(add_tc[0]), .A2(sub_tc[1]), .B(n642), .ZN(N126) );
  AOI21D0 U239 ( .A1(sub_tc[4]), .A2(n927), .B(n912), .ZN(N129) );
  OA21D0 U240 ( .A1(n639), .A2(n867), .B(n638), .Z(N132) );
  INVD0 U241 ( .I(n1210), .ZN(prod_full[23]) );
  OA21D0 U242 ( .A1(n868), .A2(n910), .B(n877), .Z(N87) );
  INVD0 U243 ( .I(n1258), .ZN(prod_full[29]) );
  INVD0 U244 ( .I(n1222), .ZN(prod_full[32]) );
  INVD0 U245 ( .I(n1182), .ZN(prod_full[35]) );
  INVD0 U246 ( .I(\mult_x_13/n207 ), .ZN(n314) );
  INVD0 U247 ( .I(\mult_x_13/n233 ), .ZN(n332) );
  INVD0 U248 ( .I(\mult_x_13/n276 ), .ZN(n350) );
  OAI22D0 U249 ( .A1(n259), .A2(n2089), .B1(n2185), .B2(n258), .ZN(n260) );
  CKND2D0 U250 ( .A1(n246), .A2(n245), .ZN(n247) );
  INVD0 U251 ( .I(\mult_x_13/n361 ), .ZN(n400) );
  INVD0 U252 ( .I(R_lat_mag[2]), .ZN(\mult_x_13/n686 ) );
  INVD0 U253 ( .I(n1194), .ZN(prod_full[14]) );
  INVD0 U254 ( .I(n76), .ZN(n74) );
  CKND2D0 U255 ( .A1(n327), .A2(n326), .ZN(n325) );
  AOI22D0 U256 ( .A1(\mult_x_13/n251 ), .A2(\mult_x_13/n259 ), .B1(n342), .B2(
        n341), .ZN(n344) );
  CKND2D0 U257 ( .A1(n373), .A2(n372), .ZN(n371) );
  CKND2D0 U258 ( .A1(n398), .A2(n397), .ZN(n396) );
  INVD0 U259 ( .I(state[0]), .ZN(n2266) );
  ND4D0 U260 ( .A1(n74), .A2(n71), .A3(n73), .A4(n72), .ZN(result_comb[1]) );
  ND4D0 U261 ( .A1(n74), .A2(n36), .A3(n38), .A4(n37), .ZN(result_comb[12]) );
  CKAN2D0 U262 ( .A1(start), .A2(n81), .Z(result_comb_valid) );
  OAI211D0 U263 ( .A1(n309), .A2(n308), .B(n412), .C(n307), .ZN(div_mag_sat[0]) );
  OAI211D0 U264 ( .A1(\mult_x_13/n260 ), .A2(n349), .B(n412), .C(n348), .ZN(
        div_mag_sat[14]) );
  CKND2D0 U265 ( .A1(ctl_d[1]), .A2(ctl_d[0]), .ZN(n81) );
  INR4D0 U266 ( .A1(start), .B1(state[0]), .B2(state[1]), .B3(n81), .ZN(N200)
         );
  BUFFD1 U267 ( .I(N200), .Z(n2267) );
  INR2XD0 U268 ( .A1(state[1]), .B1(state[0]), .ZN(n96) );
  INVD0 U269 ( .I(R_lat_mag[5]), .ZN(\mult_x_13/n660 ) );
  INVD0 U270 ( .I(S[0]), .ZN(n1418) );
  INVD0 U271 ( .I(R[14]), .ZN(n1603) );
  INVD0 U272 ( .I(R[15]), .ZN(n760) );
  AOI22D0 U273 ( .A1(R[15]), .A2(n1603), .B1(R[14]), .B2(n760), .ZN(n428) );
  NR2D0 U274 ( .A1(n1418), .A2(n428), .ZN(\mult_x_9/n382 ) );
  INVD0 U275 ( .I(R_lat_mag[17]), .ZN(\mult_x_13/n556 ) );
  INVD0 U276 ( .I(R[8]), .ZN(n1736) );
  INVD0 U277 ( .I(R[9]), .ZN(n663) );
  AOI22D0 U278 ( .A1(R[9]), .A2(n1736), .B1(R[8]), .B2(n663), .ZN(n459) );
  NR2D0 U279 ( .A1(n1418), .A2(n459), .ZN(\mult_x_9/n418 ) );
  INVD0 U280 ( .I(R_lat_mag[11]), .ZN(\mult_x_13/n608 ) );
  INVD0 U281 ( .I(R[5]), .ZN(\mult_x_9/n660 ) );
  INVD0 U282 ( .I(R[2]), .ZN(\mult_x_9/n686 ) );
  INVD0 U283 ( .I(R[11]), .ZN(\mult_x_9/n608 ) );
  INVD0 U284 ( .I(R[17]), .ZN(\mult_x_9/n556 ) );
  ND3D0 U285 ( .A1(n5), .A2(n4), .A3(n3), .ZN(n76) );
  INVD0 U286 ( .I(inv_Q_mag[0]), .ZN(n1841) );
  INVD0 U287 ( .I(R_lat_mag[6]), .ZN(n82) );
  MUX2ND0 U288 ( .I0(R_lat_mag[6]), .I1(n82), .S(R_lat_mag[7]), .ZN(n86) );
  MUX2ND0 U289 ( .I0(\mult_x_13/n660 ), .I1(R_lat_mag[5]), .S(R_lat_mag[6]), 
        .ZN(n84) );
  INVD0 U290 ( .I(n84), .ZN(n87) );
  IND2D0 U291 ( .A1(n86), .B1(n87), .ZN(n2169) );
  INVD0 U292 ( .I(inv_Q_mag[1]), .ZN(n2174) );
  INVD0 U293 ( .I(R_lat_mag[8]), .ZN(n2180) );
  MUX2ND0 U294 ( .I0(n2180), .I1(R_lat_mag[8]), .S(R_lat_mag[7]), .ZN(n88) );
  INVD0 U295 ( .I(n88), .ZN(n83) );
  CKND2D0 U296 ( .A1(n83), .A2(n84), .ZN(n2171) );
  AOI22D0 U297 ( .A1(inv_Q_mag[0]), .A2(n2174), .B1(inv_Q_mag[1]), .B2(n1841), 
        .ZN(n1843) );
  NR2D0 U298 ( .A1(n87), .A2(n83), .ZN(n2178) );
  INVD0 U299 ( .I(n2178), .ZN(n2091) );
  OA222D0 U300 ( .A1(n1841), .A2(n2169), .B1(n2174), .B2(n2171), .C1(n1843), 
        .C2(n2091), .Z(n97) );
  CKND2D0 U301 ( .A1(n84), .A2(inv_Q_mag[0]), .ZN(n118) );
  ND3D0 U302 ( .A1(R_lat_mag[8]), .A2(n97), .A3(n118), .ZN(n157) );
  INVD0 U303 ( .I(inv_Q_mag[2]), .ZN(n2170) );
  NR2D0 U304 ( .A1(inv_Q_mag[0]), .A2(n2174), .ZN(n85) );
  MUX2ND0 U305 ( .I0(n2170), .I1(inv_Q_mag[2]), .S(n85), .ZN(n1335) );
  NR2D0 U306 ( .A1(n2174), .A2(n2169), .ZN(n90) );
  ND3D0 U307 ( .A1(n88), .A2(n87), .A3(n86), .ZN(n2173) );
  OAI22D0 U308 ( .A1(n1841), .A2(n2173), .B1(n2170), .B2(n2171), .ZN(n89) );
  AOI211D0 U309 ( .A1(n2178), .A2(n1335), .B(n90), .C(n89), .ZN(n159) );
  CKND2D0 U310 ( .A1(R_lat_mag[8]), .A2(n159), .ZN(n158) );
  NR2D0 U311 ( .A1(n157), .A2(n158), .ZN(\mult_x_13/n421 ) );
  MUX2ND0 U312 ( .I0(\mult_x_13/n686 ), .I1(R_lat_mag[2]), .S(R_lat_mag[1]), 
        .ZN(n91) );
  CKND2D0 U313 ( .A1(n91), .A2(R_lat_mag[0]), .ZN(n259) );
  INVD0 U314 ( .I(n259), .ZN(n249) );
  AOI21D0 U315 ( .A1(n1841), .A2(n2170), .B(n2174), .ZN(n108) );
  NR3D0 U316 ( .A1(R_lat_mag[1]), .A2(R_lat_mag[0]), .A3(\mult_x_13/n686 ), 
        .ZN(n255) );
  AOI22D0 U317 ( .A1(n249), .A2(n2222), .B1(n255), .B2(inv_Q_mag[12]), .ZN(n93) );
  IND2D0 U318 ( .A1(R_lat_mag[0]), .B1(R_lat_mag[1]), .ZN(n256) );
  INVD0 U319 ( .I(n256), .ZN(n250) );
  INR2D0 U320 ( .A1(R_lat_mag[0]), .B1(n91), .ZN(n251) );
  AOI22D0 U321 ( .A1(n250), .A2(inv_Q_mag[13]), .B1(n251), .B2(inv_Q_mag[14]), 
        .ZN(n92) );
  CKND2D0 U322 ( .A1(n93), .A2(n92), .ZN(n94) );
  MUX2ND0 U323 ( .I0(R_lat_mag[2]), .I1(\mult_x_13/n686 ), .S(n94), .ZN(n309)
         );
  INVD0 U324 ( .I(\mult_x_13/n385 ), .ZN(n208) );
  INVD0 U325 ( .I(\mult_x_13/n392 ), .ZN(n207) );
  INVD0 U326 ( .I(\mult_x_13/n406 ), .ZN(n194) );
  OAI21D0 U327 ( .A1(n118), .A2(n2180), .B(n97), .ZN(n95) );
  OAI31D0 U328 ( .A1(n118), .A2(n97), .A3(n2180), .B(n95), .ZN(n163) );
  INVD0 U329 ( .I(n118), .ZN(n112) );
  MUX2ND0 U330 ( .I0(\mult_x_13/n686 ), .I1(R_lat_mag[2]), .S(R_lat_mag[3]), 
        .ZN(n105) );
  INVD0 U331 ( .I(R_lat_mag[3]), .ZN(n98) );
  MUX2ND0 U332 ( .I0(R_lat_mag[3]), .I1(n98), .S(R_lat_mag[4]), .ZN(n101) );
  MUX2ND0 U333 ( .I0(\mult_x_13/n660 ), .I1(R_lat_mag[5]), .S(R_lat_mag[4]), 
        .ZN(n100) );
  ND3D0 U334 ( .A1(n99), .A2(n101), .A3(n100), .ZN(n2188) );
  INVD0 U335 ( .I(n2188), .ZN(n2256) );
  CKND2D0 U336 ( .A1(n105), .A2(n100), .ZN(n2183) );
  INVD0 U337 ( .I(n2183), .ZN(n2255) );
  AOI22D0 U338 ( .A1(inv_Q_mag[0]), .A2(n2256), .B1(n1335), .B2(n2255), .ZN(
        n103) );
  NR2D0 U339 ( .A1(n100), .A2(n99), .ZN(n2258) );
  NR2D0 U340 ( .A1(n105), .A2(n101), .ZN(n2257) );
  AOI22D0 U341 ( .A1(n2258), .A2(inv_Q_mag[2]), .B1(n2257), .B2(inv_Q_mag[1]), 
        .ZN(n102) );
  CKND2D0 U342 ( .A1(n103), .A2(n102), .ZN(n104) );
  MUX2ND0 U343 ( .I0(\mult_x_13/n660 ), .I1(R_lat_mag[5]), .S(n104), .ZN(n139)
         );
  CKND2D0 U344 ( .A1(inv_Q_mag[0]), .A2(n105), .ZN(n130) );
  INR2D0 U345 ( .A1(n130), .B1(\mult_x_13/n660 ), .ZN(n107) );
  INVD0 U346 ( .I(n1843), .ZN(n557) );
  AO222D0 U347 ( .A1(inv_Q_mag[1]), .A2(n2258), .B1(n2257), .B2(inv_Q_mag[0]), 
        .C1(n2255), .C2(n557), .Z(n125) );
  INVD0 U348 ( .I(n125), .ZN(n106) );
  CKND2D0 U349 ( .A1(n107), .A2(n106), .ZN(n138) );
  INR2D0 U350 ( .A1(n139), .B1(n138), .ZN(n119) );
  FA1D0 U351 ( .A(inv_Q_mag[2]), .B(inv_Q_mag[3]), .CI(n108), .CO(n113), .S(
        n2177) );
  AOI22D0 U352 ( .A1(inv_Q_mag[1]), .A2(n2256), .B1(n2255), .B2(n2177), .ZN(
        n110) );
  AOI22D0 U353 ( .A1(n2258), .A2(inv_Q_mag[3]), .B1(inv_Q_mag[2]), .B2(n2257), 
        .ZN(n109) );
  CKND2D0 U354 ( .A1(n110), .A2(n109), .ZN(n111) );
  MUX2ND0 U355 ( .I0(\mult_x_13/n660 ), .I1(R_lat_mag[5]), .S(n111), .ZN(n117)
         );
  OAI21D0 U356 ( .A1(n112), .A2(n119), .B(n117), .ZN(n162) );
  FA1D0 U357 ( .A(inv_Q_mag[3]), .B(inv_Q_mag[4]), .CI(n113), .CO(n120), .S(
        n2167) );
  AOI22D0 U358 ( .A1(inv_Q_mag[2]), .A2(n2256), .B1(n2255), .B2(n2167), .ZN(
        n115) );
  AOI22D0 U359 ( .A1(n2258), .A2(inv_Q_mag[4]), .B1(n2257), .B2(inv_Q_mag[3]), 
        .ZN(n114) );
  CKND2D0 U360 ( .A1(n115), .A2(n114), .ZN(n116) );
  MUX2ND0 U361 ( .I0(R_lat_mag[5]), .I1(\mult_x_13/n660 ), .S(n116), .ZN(n161)
         );
  XNR3D0 U362 ( .A1(n119), .A2(n118), .A3(n117), .ZN(n149) );
  FA1D0 U363 ( .A(inv_Q_mag[4]), .B(inv_Q_mag[5]), .CI(n120), .CO(n143), .S(
        n2162) );
  AOI22D0 U364 ( .A1(n249), .A2(n2162), .B1(n255), .B2(inv_Q_mag[3]), .ZN(n122) );
  AOI22D0 U365 ( .A1(n250), .A2(inv_Q_mag[4]), .B1(n251), .B2(inv_Q_mag[5]), 
        .ZN(n121) );
  CKND2D0 U366 ( .A1(n122), .A2(n121), .ZN(n123) );
  MUX2ND0 U367 ( .I0(R_lat_mag[2]), .I1(\mult_x_13/n686 ), .S(n123), .ZN(n142)
         );
  OAI21D0 U368 ( .A1(\mult_x_13/n660 ), .A2(n130), .B(n125), .ZN(n124) );
  OAI31D0 U369 ( .A1(\mult_x_13/n660 ), .A2(n125), .A3(n130), .B(n124), .ZN(
        n137) );
  AOI22D0 U370 ( .A1(n249), .A2(n2177), .B1(n255), .B2(inv_Q_mag[1]), .ZN(n127) );
  AOI22D0 U371 ( .A1(n250), .A2(inv_Q_mag[2]), .B1(n251), .B2(inv_Q_mag[3]), 
        .ZN(n126) );
  CKND2D0 U372 ( .A1(n127), .A2(n126), .ZN(n131) );
  ND4D0 U373 ( .A1(R_lat_mag[2]), .A2(n2170), .A3(n1841), .A4(n2174), .ZN(n129) );
  NR2D0 U374 ( .A1(R_lat_mag[2]), .A2(n131), .ZN(n128) );
  AOI221D0 U375 ( .A1(R_lat_mag[2]), .A2(n131), .B1(n130), .B2(n129), .C(n128), 
        .ZN(n136) );
  AOI22D0 U376 ( .A1(n249), .A2(n2167), .B1(n255), .B2(inv_Q_mag[2]), .ZN(n133) );
  AOI22D0 U377 ( .A1(n250), .A2(inv_Q_mag[3]), .B1(n251), .B2(inv_Q_mag[4]), 
        .ZN(n132) );
  CKND2D0 U378 ( .A1(n133), .A2(n132), .ZN(n134) );
  MUX2ND0 U379 ( .I0(\mult_x_13/n686 ), .I1(R_lat_mag[2]), .S(n134), .ZN(n135)
         );
  MAOI222D0 U380 ( .A(n137), .B(n136), .C(n135), .ZN(n141) );
  CKXOR2D0 U381 ( .A1(n139), .A2(n138), .Z(n140) );
  MAOI222D0 U382 ( .A(n142), .B(n141), .C(n140), .ZN(n148) );
  FA1D0 U383 ( .A(inv_Q_mag[5]), .B(inv_Q_mag[6]), .CI(n143), .CO(n150), .S(
        n2254) );
  AOI22D0 U384 ( .A1(n249), .A2(n2254), .B1(n255), .B2(inv_Q_mag[4]), .ZN(n145) );
  AOI22D0 U385 ( .A1(n250), .A2(inv_Q_mag[5]), .B1(n251), .B2(inv_Q_mag[6]), 
        .ZN(n144) );
  CKND2D0 U386 ( .A1(n145), .A2(n144), .ZN(n146) );
  MUX2ND0 U387 ( .I0(\mult_x_13/n686 ), .I1(R_lat_mag[2]), .S(n146), .ZN(n147)
         );
  MAOI222D0 U388 ( .A(n149), .B(n148), .C(n147), .ZN(n155) );
  FA1D0 U389 ( .A(inv_Q_mag[6]), .B(inv_Q_mag[7]), .CI(n150), .CO(n168), .S(
        n2250) );
  AOI22D0 U390 ( .A1(n249), .A2(n2250), .B1(n255), .B2(inv_Q_mag[5]), .ZN(n152) );
  CKND2D0 U391 ( .A1(n152), .A2(n151), .ZN(n153) );
  MUX2ND0 U392 ( .I0(R_lat_mag[2]), .I1(\mult_x_13/n686 ), .S(n153), .ZN(n154)
         );
  MAOI222D0 U393 ( .A(n156), .B(n155), .C(n154), .ZN(n174) );
  OAI211D0 U394 ( .A1(R_lat_mag[8]), .A2(n159), .B(n158), .C(n157), .ZN(n160)
         );
  IND2D0 U395 ( .A1(\mult_x_13/n421 ), .B1(n160), .ZN(n570) );
  FA1D0 U396 ( .A(n163), .B(n162), .CI(n161), .CO(n569), .S(n156) );
  AOI22D0 U397 ( .A1(n2256), .A2(inv_Q_mag[3]), .B1(n2255), .B2(n2162), .ZN(
        n165) );
  AOI22D0 U398 ( .A1(n2258), .A2(inv_Q_mag[5]), .B1(n2257), .B2(inv_Q_mag[4]), 
        .ZN(n164) );
  CKND2D0 U399 ( .A1(n165), .A2(n164), .ZN(n166) );
  MUX2ND0 U400 ( .I0(R_lat_mag[5]), .I1(\mult_x_13/n660 ), .S(n166), .ZN(n568)
         );
  INVD0 U401 ( .I(n167), .ZN(n173) );
  FA1D0 U402 ( .A(inv_Q_mag[7]), .B(inv_Q_mag[8]), .CI(n168), .CO(n175), .S(
        n2246) );
  AOI22D0 U403 ( .A1(n249), .A2(n2246), .B1(n255), .B2(inv_Q_mag[6]), .ZN(n170) );
  AOI22D0 U404 ( .A1(n250), .A2(inv_Q_mag[7]), .B1(n251), .B2(inv_Q_mag[8]), 
        .ZN(n169) );
  MUX2ND0 U405 ( .I0(\mult_x_13/n686 ), .I1(R_lat_mag[2]), .S(n171), .ZN(n172)
         );
  MAOI222D0 U406 ( .A(n174), .B(n173), .C(n172), .ZN(n180) );
  FA1D0 U407 ( .A(inv_Q_mag[8]), .B(inv_Q_mag[9]), .CI(n175), .CO(n182), .S(
        n2242) );
  AOI22D0 U408 ( .A1(n249), .A2(n2242), .B1(n255), .B2(inv_Q_mag[7]), .ZN(n177) );
  AOI22D0 U409 ( .A1(n250), .A2(inv_Q_mag[8]), .B1(n251), .B2(inv_Q_mag[9]), 
        .ZN(n176) );
  CKND2D0 U410 ( .A1(n177), .A2(n176), .ZN(n178) );
  MUX2ND0 U411 ( .I0(R_lat_mag[2]), .I1(\mult_x_13/n686 ), .S(n178), .ZN(n179)
         );
  MAOI222D0 U412 ( .A(n181), .B(n180), .C(n179), .ZN(n187) );
  FA1D0 U413 ( .A(inv_Q_mag[9]), .B(inv_Q_mag[10]), .CI(n182), .CO(n188), .S(
        n2238) );
  AOI22D0 U414 ( .A1(n249), .A2(n2238), .B1(n255), .B2(inv_Q_mag[8]), .ZN(n184) );
  AOI22D0 U415 ( .A1(n250), .A2(inv_Q_mag[9]), .B1(n251), .B2(inv_Q_mag[10]), 
        .ZN(n183) );
  CKND2D0 U416 ( .A1(n184), .A2(n183), .ZN(n185) );
  MUX2ND0 U417 ( .I0(\mult_x_13/n686 ), .I1(R_lat_mag[2]), .S(n185), .ZN(n186)
         );
  MAOI222D0 U418 ( .A(\mult_x_13/n411 ), .B(n187), .C(n186), .ZN(n193) );
  FA1D0 U419 ( .A(inv_Q_mag[10]), .B(inv_Q_mag[11]), .CI(n188), .CO(n195), .S(
        n2234) );
  AOI22D0 U420 ( .A1(n249), .A2(n2234), .B1(n255), .B2(inv_Q_mag[9]), .ZN(n190) );
  AOI22D0 U421 ( .A1(n250), .A2(inv_Q_mag[10]), .B1(n251), .B2(inv_Q_mag[11]), 
        .ZN(n189) );
  CKND2D0 U422 ( .A1(n190), .A2(n189), .ZN(n191) );
  MUX2ND0 U423 ( .I0(R_lat_mag[2]), .I1(\mult_x_13/n686 ), .S(n191), .ZN(n192)
         );
  MAOI222D0 U424 ( .A(n194), .B(n193), .C(n192), .ZN(n200) );
  FA1D0 U425 ( .A(inv_Q_mag[11]), .B(inv_Q_mag[12]), .CI(n195), .CO(n201), .S(
        n2230) );
  AOI22D0 U426 ( .A1(n249), .A2(n2230), .B1(n255), .B2(inv_Q_mag[10]), .ZN(
        n197) );
  AOI22D0 U427 ( .A1(n250), .A2(inv_Q_mag[11]), .B1(n251), .B2(inv_Q_mag[12]), 
        .ZN(n196) );
  CKND2D0 U428 ( .A1(n197), .A2(n196), .ZN(n198) );
  MUX2ND0 U429 ( .I0(\mult_x_13/n686 ), .I1(R_lat_mag[2]), .S(n198), .ZN(n199)
         );
  MAOI222D0 U430 ( .A(\mult_x_13/n399 ), .B(n200), .C(n199), .ZN(n206) );
  FA1D0 U431 ( .A(inv_Q_mag[12]), .B(inv_Q_mag[13]), .CI(n201), .CO(n209), .S(
        n2226) );
  AOI22D0 U432 ( .A1(n249), .A2(n2226), .B1(n255), .B2(inv_Q_mag[11]), .ZN(
        n203) );
  AOI22D0 U433 ( .A1(n250), .A2(inv_Q_mag[12]), .B1(n251), .B2(inv_Q_mag[13]), 
        .ZN(n202) );
  CKND2D0 U434 ( .A1(n203), .A2(n202), .ZN(n204) );
  MUX2ND0 U435 ( .I0(R_lat_mag[2]), .I1(\mult_x_13/n686 ), .S(n204), .ZN(n205)
         );
  MAOI222D0 U436 ( .A(n207), .B(n206), .C(n205), .ZN(n220) );
  MUX2ND0 U437 ( .I0(n208), .I1(\mult_x_13/n385 ), .S(n220), .ZN(n308) );
  INVD0 U438 ( .I(R_lat_mag[20]), .ZN(n1900) );
  MUX2ND0 U439 ( .I0(n1900), .I1(R_lat_mag[20]), .S(R_lat_mag[21]), .ZN(n1380)
         );
  CKND2D0 U440 ( .A1(n1380), .A2(R_lat_mag[22]), .ZN(n1844) );
  INVD0 U441 ( .I(n1844), .ZN(n1334) );
  FA1D0 U442 ( .A(inv_Q_mag[13]), .B(inv_Q_mag[14]), .CI(n209), .CO(n221), .S(
        n2222) );
  INVD0 U443 ( .I(inv_Q_mag[18]), .ZN(n2107) );
  ND3D0 U444 ( .A1(R_lat_mag[20]), .A2(R_lat_mag[21]), .A3(R_lat_mag[22]), 
        .ZN(n1285) );
  INVD0 U445 ( .I(inv_Q_mag[20]), .ZN(n2099) );
  INVD0 U446 ( .I(R_lat_mag[22]), .ZN(n211) );
  INVD0 U447 ( .I(inv_Q_mag[19]), .ZN(n2103) );
  INVD0 U448 ( .I(R_lat_mag[21]), .ZN(n210) );
  AOI33D0 U449 ( .A1(R_lat_mag[20]), .A2(R_lat_mag[21]), .A3(n211), .B1(
        R_lat_mag[22]), .B2(n210), .B3(n1900), .ZN(n1842) );
  OAI22D0 U450 ( .A1(n2099), .A2(n1840), .B1(n2103), .B2(n1842), .ZN(n212) );
  AOI211D0 U451 ( .A1(n1334), .A2(n2198), .B(n213), .C(n212), .ZN(n268) );
  MUX2ND0 U452 ( .I0(R_lat_mag[20]), .I1(n1900), .S(R_lat_mag[19]), .ZN(n478)
         );
  MUX2ND0 U453 ( .I0(R_lat_mag[17]), .I1(\mult_x_13/n556 ), .S(R_lat_mag[18]), 
        .ZN(n479) );
  INVD0 U454 ( .I(R_lat_mag[18]), .ZN(n214) );
  MUX2ND0 U455 ( .I0(R_lat_mag[18]), .I1(n214), .S(R_lat_mag[19]), .ZN(n215)
         );
  IND3D0 U456 ( .A1(n478), .B1(n479), .B2(n215), .ZN(n1894) );
  INVD0 U457 ( .I(inv_Q_mag[21]), .ZN(n2187) );
  IND2D0 U458 ( .A1(n215), .B1(n479), .ZN(n1895) );
  INVD0 U459 ( .I(inv_Q_mag[22]), .ZN(n2185) );
  FA1D0 U460 ( .A(inv_Q_mag[19]), .B(inv_Q_mag[20]), .CI(n216), .CO(n244), .S(
        n2198) );
  OAI21D0 U461 ( .A1(inv_Q_mag[22]), .A2(n217), .B(n2089), .ZN(n2184) );
  NR2D0 U462 ( .A1(n479), .A2(n478), .ZN(n1898) );
  INVD0 U463 ( .I(n1898), .ZN(n480) );
  OAI222D0 U464 ( .A1(n1894), .A2(n2187), .B1(n1895), .B2(n2185), .C1(n2184), 
        .C2(n480), .ZN(n218) );
  MUX2ND0 U465 ( .I0(R_lat_mag[20]), .I1(n1900), .S(n218), .ZN(n267) );
  INVD0 U466 ( .I(n309), .ZN(n219) );
  MAOI222D0 U467 ( .A(\mult_x_13/n385 ), .B(n220), .C(n219), .ZN(n409) );
  FA1D0 U468 ( .A(inv_Q_mag[14]), .B(inv_Q_mag[15]), .CI(n221), .CO(n225), .S(
        n2218) );
  AOI22D0 U469 ( .A1(n249), .A2(n2218), .B1(n250), .B2(inv_Q_mag[14]), .ZN(
        n223) );
  AOI22D0 U470 ( .A1(n255), .A2(inv_Q_mag[13]), .B1(n251), .B2(inv_Q_mag[15]), 
        .ZN(n222) );
  CKND2D0 U471 ( .A1(n223), .A2(n222), .ZN(n224) );
  MUX2ND0 U472 ( .I0(R_lat_mag[2]), .I1(\mult_x_13/n686 ), .S(n224), .ZN(n414)
         );
  INVD0 U473 ( .I(\mult_x_13/n377 ), .ZN(n410) );
  MAOI222D0 U474 ( .A(n409), .B(n414), .C(n410), .ZN(n405) );
  FA1D0 U475 ( .A(inv_Q_mag[15]), .B(inv_Q_mag[16]), .CI(n225), .CO(n229), .S(
        n2214) );
  AOI22D0 U476 ( .A1(n249), .A2(n2214), .B1(n255), .B2(inv_Q_mag[14]), .ZN(
        n227) );
  AOI22D0 U477 ( .A1(n250), .A2(inv_Q_mag[15]), .B1(n251), .B2(inv_Q_mag[16]), 
        .ZN(n226) );
  CKND2D0 U478 ( .A1(n227), .A2(n226), .ZN(n228) );
  MUX2ND0 U479 ( .I0(\mult_x_13/n686 ), .I1(R_lat_mag[2]), .S(n228), .ZN(n407)
         );
  MAOI222D0 U480 ( .A(\mult_x_13/n369 ), .B(n405), .C(n407), .ZN(n399) );
  FA1D0 U481 ( .A(inv_Q_mag[16]), .B(inv_Q_mag[17]), .CI(n229), .CO(n233), .S(
        n2210) );
  AOI22D0 U482 ( .A1(n249), .A2(n2210), .B1(n255), .B2(inv_Q_mag[15]), .ZN(
        n231) );
  AOI22D0 U483 ( .A1(n250), .A2(inv_Q_mag[16]), .B1(n251), .B2(inv_Q_mag[17]), 
        .ZN(n230) );
  CKND2D0 U484 ( .A1(n231), .A2(n230), .ZN(n232) );
  MUX2ND0 U485 ( .I0(R_lat_mag[2]), .I1(\mult_x_13/n686 ), .S(n232), .ZN(n403)
         );
  MAOI222D0 U486 ( .A(n399), .B(n403), .C(n400), .ZN(n395) );
  FA1D0 U487 ( .A(inv_Q_mag[17]), .B(inv_Q_mag[18]), .CI(n233), .CO(n237), .S(
        n2206) );
  AOI22D0 U488 ( .A1(n249), .A2(n2206), .B1(n255), .B2(inv_Q_mag[16]), .ZN(
        n235) );
  AOI22D0 U489 ( .A1(n250), .A2(inv_Q_mag[17]), .B1(n251), .B2(inv_Q_mag[18]), 
        .ZN(n234) );
  CKND2D0 U490 ( .A1(n235), .A2(n234), .ZN(n236) );
  MUX2ND0 U491 ( .I0(\mult_x_13/n686 ), .I1(R_lat_mag[2]), .S(n236), .ZN(n397)
         );
  MAOI222D0 U492 ( .A(\mult_x_13/n351 ), .B(n395), .C(n397), .ZN(n389) );
  FA1D0 U493 ( .A(inv_Q_mag[18]), .B(inv_Q_mag[19]), .CI(n237), .CO(n216), .S(
        n2202) );
  AOI22D0 U494 ( .A1(n249), .A2(n2202), .B1(n255), .B2(inv_Q_mag[17]), .ZN(
        n239) );
  CKND2D0 U495 ( .A1(n239), .A2(n238), .ZN(n240) );
  MUX2ND0 U496 ( .I0(R_lat_mag[2]), .I1(\mult_x_13/n686 ), .S(n240), .ZN(n393)
         );
  INVD0 U497 ( .I(\mult_x_13/n341 ), .ZN(n390) );
  MAOI222D0 U498 ( .A(n389), .B(n393), .C(n390), .ZN(n385) );
  AOI22D0 U499 ( .A1(n249), .A2(n2198), .B1(n255), .B2(inv_Q_mag[18]), .ZN(
        n242) );
  AOI22D0 U500 ( .A1(n250), .A2(inv_Q_mag[19]), .B1(n251), .B2(inv_Q_mag[20]), 
        .ZN(n241) );
  CKND2D0 U501 ( .A1(n242), .A2(n241), .ZN(n243) );
  MUX2ND0 U502 ( .I0(\mult_x_13/n686 ), .I1(R_lat_mag[2]), .S(n243), .ZN(n387)
         );
  MAOI222D0 U503 ( .A(\mult_x_13/n331 ), .B(n385), .C(n387), .ZN(n379) );
  FA1D0 U504 ( .A(inv_Q_mag[20]), .B(inv_Q_mag[21]), .CI(n244), .CO(n248), .S(
        n2194) );
  AOI22D0 U505 ( .A1(n249), .A2(n2194), .B1(n255), .B2(inv_Q_mag[19]), .ZN(
        n246) );
  MUX2ND0 U506 ( .I0(R_lat_mag[2]), .I1(\mult_x_13/n686 ), .S(n247), .ZN(n383)
         );
  INVD0 U507 ( .I(\mult_x_13/n322 ), .ZN(n380) );
  MAOI222D0 U508 ( .A(n379), .B(n383), .C(n380), .ZN(n375) );
  FA1D0 U509 ( .A(inv_Q_mag[21]), .B(inv_Q_mag[22]), .CI(n248), .CO(n217), .S(
        n2190) );
  AOI22D0 U510 ( .A1(n249), .A2(n2190), .B1(n255), .B2(inv_Q_mag[20]), .ZN(
        n253) );
  AOI22D0 U511 ( .A1(inv_Q_mag[22]), .A2(n251), .B1(inv_Q_mag[21]), .B2(n250), 
        .ZN(n252) );
  CKND2D0 U512 ( .A1(n253), .A2(n252), .ZN(n254) );
  MUX2ND0 U513 ( .I0(\mult_x_13/n686 ), .I1(R_lat_mag[2]), .S(n254), .ZN(n377)
         );
  MAOI222D0 U514 ( .A(\mult_x_13/n313 ), .B(n375), .C(n377), .ZN(n369) );
  INVD0 U515 ( .I(n255), .ZN(n258) );
  OAI222D0 U516 ( .A1(n2187), .A2(n258), .B1(n2184), .B2(n259), .C1(n2185), 
        .C2(n256), .ZN(n257) );
  MUX2ND0 U517 ( .I0(R_lat_mag[2]), .I1(\mult_x_13/n686 ), .S(n257), .ZN(n373)
         );
  INVD0 U518 ( .I(\mult_x_13/n304 ), .ZN(n370) );
  MAOI222D0 U519 ( .A(n369), .B(n373), .C(n370), .ZN(n365) );
  MUX2ND0 U520 ( .I0(\mult_x_13/n686 ), .I1(R_lat_mag[2]), .S(n260), .ZN(n367)
         );
  MAOI222D0 U521 ( .A(\mult_x_13/n295 ), .B(n365), .C(n367), .ZN(n363) );
  INVD0 U522 ( .I(\mult_x_13/n286 ), .ZN(n359) );
  INVD0 U523 ( .I(\mult_x_13/n294 ), .ZN(n360) );
  MAOI222D0 U524 ( .A(n363), .B(n359), .C(n360), .ZN(n356) );
  MAOI222D0 U525 ( .A(\mult_x_13/n277 ), .B(\mult_x_13/n285 ), .C(n356), .ZN(
        n354) );
  INVD0 U526 ( .I(\mult_x_13/n268 ), .ZN(n351) );
  MAOI222D0 U527 ( .A(n354), .B(n350), .C(n351), .ZN(n347) );
  MAOI222D0 U528 ( .A(\mult_x_13/n260 ), .B(\mult_x_13/n267 ), .C(n347), .ZN(
        n345) );
  INVD0 U529 ( .I(\mult_x_13/n251 ), .ZN(n341) );
  INVD0 U530 ( .I(\mult_x_13/n259 ), .ZN(n342) );
  MAOI222D0 U531 ( .A(n345), .B(n341), .C(n342), .ZN(n338) );
  MAOI222D0 U532 ( .A(\mult_x_13/n250 ), .B(\mult_x_13/n241 ), .C(n338), .ZN(
        n336) );
  INVD0 U533 ( .I(\mult_x_13/n240 ), .ZN(n333) );
  MAOI222D0 U534 ( .A(n336), .B(n332), .C(n333), .ZN(n329) );
  MAOI222D0 U535 ( .A(\mult_x_13/n226 ), .B(\mult_x_13/n232 ), .C(n329), .ZN(
        n327) );
  INVD0 U536 ( .I(\mult_x_13/n225 ), .ZN(n323) );
  INVD0 U537 ( .I(\mult_x_13/n218 ), .ZN(n324) );
  MAOI222D0 U538 ( .A(n327), .B(n323), .C(n324), .ZN(n320) );
  MAOI222D0 U539 ( .A(\mult_x_13/n213 ), .B(\mult_x_13/n217 ), .C(n320), .ZN(
        n318) );
  INVD0 U540 ( .I(\mult_x_13/n212 ), .ZN(n315) );
  MAOI222D0 U541 ( .A(n318), .B(n314), .C(n315), .ZN(n311) );
  MAOI222D0 U542 ( .A(\mult_x_13/n206 ), .B(\mult_x_13/n200 ), .C(n311), .ZN(
        n287) );
  INVD0 U543 ( .I(\mult_x_13/n196 ), .ZN(n281) );
  CKND2D0 U544 ( .A1(n287), .A2(n281), .ZN(n277) );
  NR2D0 U545 ( .A1(\mult_x_13/n192 ), .A2(n277), .ZN(n284) );
  CKND2D0 U546 ( .A1(n284), .A2(n282), .ZN(n288) );
  NR2D0 U547 ( .A1(\mult_x_13/n184 ), .A2(n288), .ZN(n261) );
  OAI22D0 U548 ( .A1(n2185), .A2(n1894), .B1(n2089), .B2(n480), .ZN(n263) );
  MUX2ND0 U549 ( .I0(R_lat_mag[20]), .I1(n1900), .S(n263), .ZN(n291) );
  NR2D0 U550 ( .A1(n2103), .A2(n1285), .ZN(n265) );
  OAI22D0 U551 ( .A1(n2187), .A2(n1840), .B1(n2099), .B2(n1842), .ZN(n264) );
  AOI211D0 U552 ( .A1(n1334), .A2(n2194), .B(n265), .C(n264), .ZN(n290) );
  INVD0 U553 ( .I(n273), .ZN(n266) );
  MUX2ND0 U554 ( .I0(n273), .I1(n266), .S(n274), .ZN(n271) );
  FA1D0 U555 ( .A(\mult_x_13/n178 ), .B(n268), .CI(n267), .CO(n270), .S(n262)
         );
  OAI22D0 U556 ( .A1(\mult_x_13/n183 ), .A2(n272), .B1(n271), .B2(n270), .ZN(
        n269) );
  AOI221D0 U557 ( .A1(n272), .A2(\mult_x_13/n183 ), .B1(n271), .B2(n270), .C(
        n269), .ZN(n306) );
  IND2D0 U558 ( .A1(n274), .B1(n273), .ZN(n293) );
  OAI222D0 U559 ( .A1(n1285), .A2(n2187), .B1(n1842), .B2(n2185), .C1(n1844), 
        .C2(n2184), .ZN(n279) );
  NR2D0 U560 ( .A1(n2099), .A2(n1285), .ZN(n276) );
  OAI22D0 U561 ( .A1(n2185), .A2(n1840), .B1(n2187), .B2(n1842), .ZN(n275) );
  AO211D0 U562 ( .A1(n1334), .A2(n2190), .B(n276), .C(n275), .Z(n292) );
  OA21D0 U563 ( .A1(n1900), .A2(\mult_x_13/n178 ), .B(n292), .Z(n278) );
  INVD0 U564 ( .I(n1285), .ZN(n1337) );
  AOI22D0 U565 ( .A1(inv_Q_mag[22]), .A2(n1337), .B1(n2181), .B2(n1334), .ZN(
        n280) );
  AOI31D0 U566 ( .A1(n293), .A2(n279), .A3(n278), .B(n280), .ZN(n305) );
  XOR3D0 U567 ( .A1(\mult_x_13/n192 ), .A2(n277), .A3(\mult_x_13/n195 ), .Z(
        n304) );
  NR2D0 U568 ( .A1(n279), .A2(n278), .ZN(n302) );
  MUX2ND0 U569 ( .I0(n281), .I1(\mult_x_13/n196 ), .S(\mult_x_13/n199 ), .ZN(
        n286) );
  MUX2ND0 U570 ( .I0(n282), .I1(\mult_x_13/n191 ), .S(\mult_x_13/n187 ), .ZN(
        n285) );
  OAI22D0 U571 ( .A1(n287), .A2(n286), .B1(n284), .B2(n285), .ZN(n283) );
  AOI221D0 U572 ( .A1(n287), .A2(n286), .B1(n285), .B2(n284), .C(n283), .ZN(
        n300) );
  INVD0 U573 ( .I(\mult_x_13/n184 ), .ZN(n289) );
  MUX2ND0 U574 ( .I0(n289), .I1(\mult_x_13/n184 ), .S(\mult_x_13/n186 ), .ZN(
        n297) );
  FA1D0 U575 ( .A(\mult_x_13/n178 ), .B(n291), .CI(n290), .CO(n294), .S(n273)
         );
  XNR4D0 U576 ( .A1(\mult_x_13/n178 ), .A2(n294), .A3(n293), .A4(n292), .ZN(
        n296) );
  OAI22D0 U577 ( .A1(n298), .A2(n297), .B1(n296), .B2(R_lat_mag[20]), .ZN(n295) );
  AOI221D0 U578 ( .A1(n298), .A2(n297), .B1(R_lat_mag[20]), .B2(n296), .C(n295), .ZN(n299) );
  OAI211D0 U579 ( .A1(n302), .A2(n301), .B(n300), .C(n299), .ZN(n303) );
  INR4D0 U580 ( .A1(n306), .B1(n305), .B2(n304), .B3(n303), .ZN(n412) );
  CKND2D0 U581 ( .A1(n309), .A2(n308), .ZN(n307) );
  INVD0 U582 ( .I(n311), .ZN(n310) );
  MUX2ND0 U583 ( .I0(n311), .I1(n310), .S(\mult_x_13/n200 ), .ZN(n313) );
  CKND2D0 U584 ( .A1(\mult_x_13/n206 ), .A2(n313), .ZN(n312) );
  OAI211D0 U585 ( .A1(\mult_x_13/n206 ), .A2(n313), .B(n412), .C(n312), .ZN(
        div_mag_sat[22]) );
  AOI22D0 U586 ( .A1(\mult_x_13/n207 ), .A2(\mult_x_13/n212 ), .B1(n315), .B2(
        n314), .ZN(n317) );
  CKND2D0 U587 ( .A1(n318), .A2(n317), .ZN(n316) );
  OAI211D0 U588 ( .A1(n318), .A2(n317), .B(n412), .C(n316), .ZN(
        div_mag_sat[21]) );
  INVD0 U589 ( .I(n320), .ZN(n319) );
  MUX2ND0 U590 ( .I0(n320), .I1(n319), .S(\mult_x_13/n217 ), .ZN(n322) );
  CKND2D0 U591 ( .A1(\mult_x_13/n213 ), .A2(n322), .ZN(n321) );
  OAI211D0 U592 ( .A1(\mult_x_13/n213 ), .A2(n322), .B(n412), .C(n321), .ZN(
        div_mag_sat[20]) );
  AOI22D0 U593 ( .A1(\mult_x_13/n225 ), .A2(\mult_x_13/n218 ), .B1(n324), .B2(
        n323), .ZN(n326) );
  OAI211D0 U594 ( .A1(n327), .A2(n326), .B(n412), .C(n325), .ZN(
        div_mag_sat[19]) );
  INVD0 U595 ( .I(n329), .ZN(n328) );
  MUX2ND0 U596 ( .I0(n329), .I1(n328), .S(\mult_x_13/n232 ), .ZN(n331) );
  CKND2D0 U597 ( .A1(\mult_x_13/n226 ), .A2(n331), .ZN(n330) );
  OAI211D0 U598 ( .A1(\mult_x_13/n226 ), .A2(n331), .B(n412), .C(n330), .ZN(
        div_mag_sat[18]) );
  AOI22D0 U599 ( .A1(\mult_x_13/n233 ), .A2(\mult_x_13/n240 ), .B1(n333), .B2(
        n332), .ZN(n335) );
  CKND2D0 U600 ( .A1(n336), .A2(n335), .ZN(n334) );
  OAI211D0 U601 ( .A1(n336), .A2(n335), .B(n412), .C(n334), .ZN(
        div_mag_sat[17]) );
  INVD0 U602 ( .I(n338), .ZN(n337) );
  MUX2ND0 U603 ( .I0(n338), .I1(n337), .S(\mult_x_13/n241 ), .ZN(n340) );
  CKND2D0 U604 ( .A1(\mult_x_13/n250 ), .A2(n340), .ZN(n339) );
  OAI211D0 U605 ( .A1(\mult_x_13/n250 ), .A2(n340), .B(n412), .C(n339), .ZN(
        div_mag_sat[16]) );
  CKND2D0 U606 ( .A1(n345), .A2(n344), .ZN(n343) );
  OAI211D0 U607 ( .A1(n345), .A2(n344), .B(n412), .C(n343), .ZN(
        div_mag_sat[15]) );
  INVD0 U608 ( .I(n347), .ZN(n346) );
  MUX2ND0 U609 ( .I0(n347), .I1(n346), .S(\mult_x_13/n267 ), .ZN(n349) );
  CKND2D0 U610 ( .A1(\mult_x_13/n260 ), .A2(n349), .ZN(n348) );
  AOI22D0 U611 ( .A1(\mult_x_13/n276 ), .A2(\mult_x_13/n268 ), .B1(n351), .B2(
        n350), .ZN(n353) );
  CKND2D0 U612 ( .A1(n354), .A2(n353), .ZN(n352) );
  OAI211D0 U613 ( .A1(n354), .A2(n353), .B(n412), .C(n352), .ZN(
        div_mag_sat[13]) );
  INVD0 U614 ( .I(n356), .ZN(n355) );
  MUX2ND0 U615 ( .I0(n356), .I1(n355), .S(\mult_x_13/n285 ), .ZN(n358) );
  CKND2D0 U616 ( .A1(\mult_x_13/n277 ), .A2(n358), .ZN(n357) );
  OAI211D0 U617 ( .A1(\mult_x_13/n277 ), .A2(n358), .B(n412), .C(n357), .ZN(
        div_mag_sat[12]) );
  AOI22D0 U618 ( .A1(\mult_x_13/n286 ), .A2(\mult_x_13/n294 ), .B1(n360), .B2(
        n359), .ZN(n362) );
  CKND2D0 U619 ( .A1(n363), .A2(n362), .ZN(n361) );
  OAI211D0 U620 ( .A1(n363), .A2(n362), .B(n412), .C(n361), .ZN(
        div_mag_sat[11]) );
  INVD0 U621 ( .I(n365), .ZN(n364) );
  MUX2ND0 U622 ( .I0(n365), .I1(n364), .S(\mult_x_13/n295 ), .ZN(n368) );
  CKND2D0 U623 ( .A1(n368), .A2(n367), .ZN(n366) );
  OAI211D0 U624 ( .A1(n368), .A2(n367), .B(n412), .C(n366), .ZN(
        div_mag_sat[10]) );
  MUX2ND0 U625 ( .I0(\mult_x_13/n304 ), .I1(n370), .S(n369), .ZN(n372) );
  OAI211D0 U626 ( .A1(n373), .A2(n372), .B(n412), .C(n371), .ZN(div_mag_sat[9]) );
  INVD0 U627 ( .I(n375), .ZN(n374) );
  MUX2ND0 U628 ( .I0(n375), .I1(n374), .S(\mult_x_13/n313 ), .ZN(n378) );
  CKND2D0 U629 ( .A1(n378), .A2(n377), .ZN(n376) );
  OAI211D0 U630 ( .A1(n378), .A2(n377), .B(n412), .C(n376), .ZN(div_mag_sat[8]) );
  MUX2ND0 U631 ( .I0(\mult_x_13/n322 ), .I1(n380), .S(n379), .ZN(n382) );
  CKND2D0 U632 ( .A1(n383), .A2(n382), .ZN(n381) );
  OAI211D0 U633 ( .A1(n383), .A2(n382), .B(n412), .C(n381), .ZN(div_mag_sat[7]) );
  INVD0 U634 ( .I(n385), .ZN(n384) );
  MUX2ND0 U635 ( .I0(n385), .I1(n384), .S(\mult_x_13/n331 ), .ZN(n388) );
  CKND2D0 U636 ( .A1(n388), .A2(n387), .ZN(n386) );
  OAI211D0 U637 ( .A1(n388), .A2(n387), .B(n412), .C(n386), .ZN(div_mag_sat[6]) );
  MUX2ND0 U638 ( .I0(\mult_x_13/n341 ), .I1(n390), .S(n389), .ZN(n392) );
  CKND2D0 U639 ( .A1(n393), .A2(n392), .ZN(n391) );
  OAI211D0 U640 ( .A1(n393), .A2(n392), .B(n412), .C(n391), .ZN(div_mag_sat[5]) );
  INVD0 U641 ( .I(n395), .ZN(n394) );
  MUX2ND0 U642 ( .I0(n395), .I1(n394), .S(\mult_x_13/n351 ), .ZN(n398) );
  OAI211D0 U643 ( .A1(n398), .A2(n397), .B(n412), .C(n396), .ZN(div_mag_sat[4]) );
  MUX2ND0 U644 ( .I0(\mult_x_13/n361 ), .I1(n400), .S(n399), .ZN(n402) );
  CKND2D0 U645 ( .A1(n403), .A2(n402), .ZN(n401) );
  OAI211D0 U646 ( .A1(n403), .A2(n402), .B(n412), .C(n401), .ZN(div_mag_sat[3]) );
  INVD0 U647 ( .I(n405), .ZN(n404) );
  MUX2ND0 U648 ( .I0(n405), .I1(n404), .S(\mult_x_13/n369 ), .ZN(n408) );
  CKND2D0 U649 ( .A1(n408), .A2(n407), .ZN(n406) );
  OAI211D0 U650 ( .A1(n408), .A2(n407), .B(n412), .C(n406), .ZN(div_mag_sat[2]) );
  MUX2ND0 U651 ( .I0(\mult_x_13/n377 ), .I1(n410), .S(n409), .ZN(n413) );
  CKND2D0 U652 ( .A1(n414), .A2(n413), .ZN(n411) );
  OAI211D0 U653 ( .A1(n414), .A2(n413), .B(n412), .C(n411), .ZN(div_mag_sat[1]) );
  IND2D0 U654 ( .A1(done), .B1(N200), .ZN(n415) );
  INVD0 U655 ( .I(n415), .ZN(inv_start) );
  OAI31D0 U656 ( .A1(state[1]), .A2(inv_rdy), .A3(n2266), .B(n415), .ZN(
        next_state[0]) );
  INVD0 U657 ( .I(R[18]), .ZN(n744) );
  AOI22D0 U658 ( .A1(R[18]), .A2(\mult_x_9/n556 ), .B1(R[17]), .B2(n744), .ZN(
        n418) );
  NR2D0 U659 ( .A1(n1418), .A2(n418), .ZN(n1400) );
  INVD0 U660 ( .I(R[20]), .ZN(n1477) );
  INVD0 U661 ( .I(R[19]), .ZN(n765) );
  AOI22D0 U662 ( .A1(R[20]), .A2(R[19]), .B1(n765), .B2(n1477), .ZN(n419) );
  INR2D0 U663 ( .A1(n419), .B1(n418), .ZN(n1475) );
  INVD0 U664 ( .I(S[1]), .ZN(n1728) );
  CKND2D0 U665 ( .A1(n1418), .A2(n1728), .ZN(n601) );
  CKND2D0 U666 ( .A1(S[0]), .A2(S[1]), .ZN(n416) );
  CKND2D0 U667 ( .A1(n601), .A2(n416), .ZN(n1420) );
  OAI22D0 U668 ( .A1(n765), .A2(n744), .B1(R[18]), .B2(R[19]), .ZN(n417) );
  IND2D0 U669 ( .A1(n417), .B1(n418), .ZN(n1472) );
  NR2D0 U670 ( .A1(n418), .A2(n419), .ZN(n423) );
  INVD0 U671 ( .I(n423), .ZN(n1470) );
  OAI222D0 U672 ( .A1(n1037), .A2(n1420), .B1(n1472), .B2(n1418), .C1(n1470), 
        .C2(n1728), .ZN(n442) );
  OR3D0 U673 ( .A1(n1400), .A2(n1477), .A3(n442), .Z(n424) );
  NR2D0 U674 ( .A1(n1728), .A2(n1472), .ZN(n422) );
  ND3D0 U675 ( .A1(n419), .A2(n418), .A3(n417), .ZN(n1471) );
  INVD0 U676 ( .I(S[2]), .ZN(n1726) );
  NR2D0 U677 ( .A1(S[0]), .A2(n1728), .ZN(n420) );
  MUX2ND0 U678 ( .I0(S[2]), .I1(n1726), .S(n420), .ZN(n1325) );
  OAI22D0 U679 ( .A1(n1418), .A2(n1471), .B1(n1325), .B2(n1037), .ZN(n421) );
  AOI211D0 U680 ( .A1(n423), .A2(S[2]), .B(n422), .C(n421), .ZN(n426) );
  NR2D0 U681 ( .A1(n424), .A2(n425), .ZN(\mult_x_9/n337 ) );
  OAI211D0 U682 ( .A1(R[20]), .A2(n426), .B(n425), .C(n424), .ZN(n427) );
  IND2D0 U683 ( .A1(\mult_x_9/n337 ), .B1(n427), .ZN(n1342) );
  INVD0 U684 ( .I(R[16]), .ZN(n751) );
  OAI22D0 U685 ( .A1(\mult_x_9/n556 ), .A2(n751), .B1(R[16]), .B2(R[17]), .ZN(
        n429) );
  NR2D0 U686 ( .A1(n428), .A2(n429), .ZN(n1534) );
  AOI21D0 U687 ( .A1(n1726), .A2(n1418), .B(n1728), .ZN(n437) );
  INVD0 U688 ( .I(S[4]), .ZN(n1825) );
  INVD0 U689 ( .I(n428), .ZN(n431) );
  CKND2D0 U690 ( .A1(n429), .A2(n431), .ZN(n1529) );
  NR2D0 U691 ( .A1(n1825), .A2(n1529), .ZN(n433) );
  INVD0 U692 ( .I(S[3]), .ZN(n1730) );
  AOI22D0 U693 ( .A1(R[16]), .A2(R[15]), .B1(n760), .B2(n751), .ZN(n430) );
  CKND2D0 U694 ( .A1(n428), .A2(n430), .ZN(n1531) );
  OR3D0 U695 ( .A1(n431), .A2(n430), .A3(n429), .Z(n1530) );
  OAI22D0 U696 ( .A1(n1730), .A2(n1531), .B1(n1726), .B2(n1530), .ZN(n432) );
  AOI211D0 U697 ( .A1(n1534), .A2(n1723), .B(n433), .C(n432), .ZN(n434) );
  MUX2ND0 U698 ( .I0(\mult_x_9/n556 ), .I1(R[17]), .S(n434), .ZN(n1328) );
  INVD0 U699 ( .I(n1534), .ZN(n1479) );
  OA22D0 U700 ( .A1(n1418), .A2(n1530), .B1(n1728), .B2(n1531), .Z(n436) );
  OR2D0 U701 ( .A1(n1529), .A2(n1726), .Z(n435) );
  OAI211D0 U702 ( .A1(n1325), .A2(n1479), .B(n436), .C(n435), .ZN(n1316) );
  NR2D0 U703 ( .A1(\mult_x_9/n556 ), .A2(n1316), .ZN(n1314) );
  OAI222D0 U704 ( .A1(n1479), .A2(n1420), .B1(n1531), .B2(n1418), .C1(n1728), 
        .C2(n1529), .ZN(n1413) );
  NR3D0 U705 ( .A1(\mult_x_9/n382 ), .A2(\mult_x_9/n556 ), .A3(n1413), .ZN(
        n1315) );
  CKAN2D0 U706 ( .A1(n1314), .A2(n1315), .Z(n1399) );
  FA1D0 U707 ( .A(S[2]), .B(S[3]), .CI(n437), .CO(n444), .S(n1733) );
  NR2D0 U708 ( .A1(n1730), .A2(n1529), .ZN(n439) );
  OAI22D0 U709 ( .A1(n1726), .A2(n1531), .B1(n1728), .B2(n1530), .ZN(n438) );
  AOI211D0 U710 ( .A1(n1534), .A2(n1733), .B(n439), .C(n438), .ZN(n440) );
  MUX2ND0 U711 ( .I0(R[17]), .I1(\mult_x_9/n556 ), .S(n440), .ZN(n1398) );
  OAI21D0 U712 ( .A1(n1399), .A2(n1400), .B(n1398), .ZN(n1327) );
  INVD0 U713 ( .I(n442), .ZN(n443) );
  CKND2D0 U714 ( .A1(R[20]), .A2(n1400), .ZN(n441) );
  MUX2ND0 U715 ( .I0(n443), .I1(n442), .S(n441), .ZN(n1326) );
  FA1D0 U716 ( .A(S[3]), .B(S[4]), .CI(n444), .CO(n572), .S(n1723) );
  INVD0 U717 ( .I(S[5]), .ZN(n1827) );
  NR2D0 U718 ( .A1(n1827), .A2(n1529), .ZN(n446) );
  OAI22D0 U719 ( .A1(n1825), .A2(n1531), .B1(n1730), .B2(n1530), .ZN(n445) );
  AOI211D0 U720 ( .A1(n1534), .A2(n1719), .B(n446), .C(n445), .ZN(n447) );
  MUX2ND0 U721 ( .I0(\mult_x_9/n556 ), .I1(R[17]), .S(n447), .ZN(n1340) );
  INVD0 U722 ( .I(n448), .ZN(\mult_x_9/n335 ) );
  INVD0 U723 ( .I(R[12]), .ZN(n693) );
  AOI22D0 U724 ( .A1(R[12]), .A2(\mult_x_9/n608 ), .B1(R[11]), .B2(n693), .ZN(
        n450) );
  NR2D0 U725 ( .A1(n1418), .A2(n450), .ZN(n1406) );
  INVD0 U726 ( .I(R[13]), .ZN(n711) );
  AOI22D0 U727 ( .A1(R[14]), .A2(R[13]), .B1(n711), .B2(n1603), .ZN(n451) );
  INR2D0 U728 ( .A1(n451), .B1(n450), .ZN(n1601) );
  OAI22D0 U729 ( .A1(n711), .A2(n693), .B1(R[12]), .B2(R[13]), .ZN(n449) );
  IND2D0 U730 ( .A1(n449), .B1(n450), .ZN(n1596) );
  NR2D0 U731 ( .A1(n450), .A2(n451), .ZN(n454) );
  INVD0 U732 ( .I(n454), .ZN(n1598) );
  OAI222D0 U733 ( .A1(n1537), .A2(n1420), .B1(n1596), .B2(n1418), .C1(n1728), 
        .C2(n1598), .ZN(n472) );
  OR3D0 U734 ( .A1(n1406), .A2(n1603), .A3(n472), .Z(n455) );
  NR2D0 U735 ( .A1(n1728), .A2(n1596), .ZN(n453) );
  ND3D0 U736 ( .A1(n451), .A2(n450), .A3(n449), .ZN(n1597) );
  OAI22D0 U737 ( .A1(n1418), .A2(n1597), .B1(n1325), .B2(n1537), .ZN(n452) );
  AOI211D0 U738 ( .A1(n454), .A2(S[2]), .B(n453), .C(n452), .ZN(n457) );
  CKND2D0 U739 ( .A1(R[14]), .A2(n457), .ZN(n456) );
  NR2D0 U740 ( .A1(n455), .A2(n456), .ZN(\mult_x_9/n388 ) );
  OAI211D0 U741 ( .A1(R[14]), .A2(n457), .B(n456), .C(n455), .ZN(n458) );
  IND2D0 U742 ( .A1(\mult_x_9/n388 ), .B1(n458), .ZN(n1350) );
  INVD0 U743 ( .I(R[10]), .ZN(n700) );
  OAI22D0 U744 ( .A1(\mult_x_9/n608 ), .A2(n700), .B1(R[10]), .B2(R[11]), .ZN(
        n460) );
  NR2D0 U745 ( .A1(n459), .A2(n460), .ZN(n1660) );
  INVD0 U746 ( .I(n459), .ZN(n462) );
  CKND2D0 U747 ( .A1(n460), .A2(n462), .ZN(n1655) );
  NR2D0 U748 ( .A1(n1825), .A2(n1655), .ZN(n464) );
  AOI22D0 U749 ( .A1(R[10]), .A2(R[9]), .B1(n663), .B2(n700), .ZN(n461) );
  CKND2D0 U750 ( .A1(n459), .A2(n461), .ZN(n1657) );
  OR3D0 U751 ( .A1(n462), .A2(n461), .A3(n460), .Z(n1656) );
  OAI22D0 U752 ( .A1(n1730), .A2(n1657), .B1(n1726), .B2(n1656), .ZN(n463) );
  AOI211D0 U753 ( .A1(n1660), .A2(n1723), .B(n464), .C(n463), .ZN(n465) );
  MUX2ND0 U754 ( .I0(\mult_x_9/n608 ), .I1(R[11]), .S(n465), .ZN(n1358) );
  INVD0 U755 ( .I(n1660), .ZN(n1605) );
  OA22D0 U756 ( .A1(n1418), .A2(n1656), .B1(n1728), .B2(n1657), .Z(n467) );
  OR2D0 U757 ( .A1(n1655), .A2(n1726), .Z(n466) );
  OAI211D0 U758 ( .A1(n1325), .A2(n1605), .B(n467), .C(n466), .ZN(n1354) );
  NR2D0 U759 ( .A1(\mult_x_9/n608 ), .A2(n1354), .ZN(n1352) );
  OAI222D0 U760 ( .A1(n1605), .A2(n1420), .B1(n1657), .B2(n1418), .C1(n1728), 
        .C2(n1655), .ZN(n1416) );
  NR3D0 U761 ( .A1(\mult_x_9/n418 ), .A2(\mult_x_9/n608 ), .A3(n1416), .ZN(
        n1353) );
  CKAN2D0 U762 ( .A1(n1352), .A2(n1353), .Z(n1405) );
  NR2D0 U763 ( .A1(n1730), .A2(n1655), .ZN(n469) );
  OAI22D0 U764 ( .A1(n1726), .A2(n1657), .B1(n1728), .B2(n1656), .ZN(n468) );
  AOI211D0 U765 ( .A1(n1660), .A2(n1733), .B(n469), .C(n468), .ZN(n470) );
  MUX2ND0 U766 ( .I0(R[11]), .I1(\mult_x_9/n608 ), .S(n470), .ZN(n1404) );
  OAI21D0 U767 ( .A1(n1405), .A2(n1406), .B(n1404), .ZN(n1357) );
  INVD0 U768 ( .I(n472), .ZN(n473) );
  CKND2D0 U769 ( .A1(R[14]), .A2(n1406), .ZN(n471) );
  MUX2ND0 U770 ( .I0(n473), .I1(n472), .S(n471), .ZN(n1356) );
  NR2D0 U771 ( .A1(n1827), .A2(n1655), .ZN(n475) );
  MUX2ND0 U772 ( .I0(\mult_x_9/n608 ), .I1(R[11]), .S(n476), .ZN(n1348) );
  INVD0 U773 ( .I(n477), .ZN(\mult_x_9/n386 ) );
  NR2D0 U774 ( .A1(n1841), .A2(n479), .ZN(n1403) );
  IND2D0 U775 ( .A1(n479), .B1(n478), .ZN(n1893) );
  OAI222D0 U776 ( .A1(n480), .A2(n1843), .B1(n1895), .B2(n1841), .C1(n1893), 
        .C2(n2174), .ZN(n501) );
  OR3D0 U777 ( .A1(n1403), .A2(n1900), .A3(n501), .Z(n483) );
  NR2D0 U778 ( .A1(n2170), .A2(n1893), .ZN(n482) );
  OAI22D0 U779 ( .A1(n1841), .A2(n1894), .B1(n2174), .B2(n1895), .ZN(n481) );
  AOI211D0 U780 ( .A1(n1898), .A2(n1335), .B(n482), .C(n481), .ZN(n485) );
  CKND2D0 U781 ( .A1(R_lat_mag[20]), .A2(n485), .ZN(n484) );
  NR2D0 U782 ( .A1(n483), .A2(n484), .ZN(\mult_x_13/n337 ) );
  INVD0 U783 ( .I(R_lat_mag[14]), .ZN(n2028) );
  MUX2ND0 U784 ( .I0(R_lat_mag[14]), .I1(n2028), .S(R_lat_mag[15]), .ZN(n490)
         );
  NR2D0 U785 ( .A1(n1841), .A2(n490), .ZN(\mult_x_13/n382 ) );
  OAI211D0 U786 ( .A1(R_lat_mag[20]), .A2(n485), .B(n484), .C(n483), .ZN(n486)
         );
  IND2D0 U787 ( .A1(\mult_x_13/n337 ), .B1(n486), .ZN(n1346) );
  INVD0 U788 ( .I(R_lat_mag[15]), .ZN(n487) );
  MUX2ND0 U789 ( .I0(R_lat_mag[15]), .I1(n487), .S(R_lat_mag[16]), .ZN(n488)
         );
  MUX2ND0 U790 ( .I0(\mult_x_13/n556 ), .I1(R_lat_mag[17]), .S(R_lat_mag[16]), 
        .ZN(n491) );
  ND3D0 U791 ( .A1(n490), .A2(n488), .A3(n491), .ZN(n1904) );
  INVD0 U792 ( .I(n1904), .ZN(n1955) );
  INVD0 U793 ( .I(n490), .ZN(n489) );
  CKND2D0 U794 ( .A1(n489), .A2(n491), .ZN(n1902) );
  INVD0 U795 ( .I(n1902), .ZN(n1954) );
  AOI22D0 U796 ( .A1(inv_Q_mag[2]), .A2(n1955), .B1(n2167), .B2(n1954), .ZN(
        n493) );
  NR2D0 U797 ( .A1(n489), .A2(n488), .ZN(n1957) );
  NR2D0 U798 ( .A1(n491), .A2(n490), .ZN(n1956) );
  AOI22D0 U799 ( .A1(inv_Q_mag[3]), .A2(n1957), .B1(inv_Q_mag[4]), .B2(n1956), 
        .ZN(n492) );
  CKND2D0 U800 ( .A1(n493), .A2(n492), .ZN(n494) );
  MUX2ND0 U801 ( .I0(R_lat_mag[17]), .I1(\mult_x_13/n556 ), .S(n494), .ZN(
        n1332) );
  AOI22D0 U802 ( .A1(inv_Q_mag[0]), .A2(n1955), .B1(n1335), .B2(n1954), .ZN(
        n496) );
  AOI22D0 U803 ( .A1(inv_Q_mag[2]), .A2(n1956), .B1(inv_Q_mag[1]), .B2(n1957), 
        .ZN(n495) );
  CKND2D0 U804 ( .A1(n496), .A2(n495), .ZN(n1320) );
  NR2D0 U805 ( .A1(\mult_x_13/n556 ), .A2(n1320), .ZN(n1318) );
  AOI222D0 U806 ( .A1(n1954), .A2(n557), .B1(n1957), .B2(inv_Q_mag[0]), .C1(
        inv_Q_mag[1]), .C2(n1956), .ZN(n1835) );
  INVD0 U807 ( .I(n1835), .ZN(n1836) );
  NR3D0 U808 ( .A1(\mult_x_13/n382 ), .A2(\mult_x_13/n556 ), .A3(n1836), .ZN(
        n1319) );
  CKAN2D0 U809 ( .A1(n1318), .A2(n1319), .Z(n1402) );
  AOI22D0 U810 ( .A1(inv_Q_mag[1]), .A2(n1955), .B1(n2177), .B2(n1954), .ZN(
        n498) );
  AOI22D0 U811 ( .A1(inv_Q_mag[2]), .A2(n1957), .B1(inv_Q_mag[3]), .B2(n1956), 
        .ZN(n497) );
  CKND2D0 U812 ( .A1(n498), .A2(n497), .ZN(n499) );
  MUX2ND0 U813 ( .I0(\mult_x_13/n556 ), .I1(R_lat_mag[17]), .S(n499), .ZN(
        n1401) );
  OAI21D0 U814 ( .A1(n1402), .A2(n1403), .B(n1401), .ZN(n1331) );
  INVD0 U815 ( .I(n501), .ZN(n502) );
  CKND2D0 U816 ( .A1(R_lat_mag[20]), .A2(n1403), .ZN(n500) );
  MUX2ND0 U817 ( .I0(n502), .I1(n501), .S(n500), .ZN(n1330) );
  AOI22D0 U818 ( .A1(inv_Q_mag[3]), .A2(n1955), .B1(n2162), .B2(n1954), .ZN(
        n504) );
  CKND2D0 U819 ( .A1(n504), .A2(n503), .ZN(n505) );
  MUX2ND0 U820 ( .I0(R_lat_mag[17]), .I1(\mult_x_13/n556 ), .S(n505), .ZN(
        n1344) );
  INVD0 U821 ( .I(n506), .ZN(\mult_x_13/n335 ) );
  INVD0 U822 ( .I(R[6]), .ZN(n589) );
  AOI22D0 U823 ( .A1(R[6]), .A2(R[5]), .B1(\mult_x_9/n660 ), .B2(n589), .ZN(
        n513) );
  INVD0 U824 ( .I(R[7]), .ZN(n612) );
  AOI22D0 U825 ( .A1(R[7]), .A2(R[6]), .B1(n589), .B2(n612), .ZN(n507) );
  AOI22D0 U826 ( .A1(R[8]), .A2(n612), .B1(R[7]), .B2(n1736), .ZN(n508) );
  NR3D0 U827 ( .A1(n513), .A2(n507), .A3(n508), .ZN(n1662) );
  INVD0 U828 ( .I(n513), .ZN(n509) );
  CKND2D0 U829 ( .A1(n507), .A2(n509), .ZN(n1725) );
  NR2D0 U830 ( .A1(n1728), .A2(n1725), .ZN(n511) );
  CKND2D0 U831 ( .A1(n513), .A2(n508), .ZN(n1729) );
  NR2D0 U832 ( .A1(n509), .A2(n508), .ZN(n1734) );
  INVD0 U833 ( .I(n1734), .ZN(n1664) );
  OAI22D0 U834 ( .A1(n1726), .A2(n1729), .B1(n1325), .B2(n1664), .ZN(n510) );
  AOI211D0 U835 ( .A1(S[0]), .A2(n1662), .B(n511), .C(n510), .ZN(n512) );
  MUX2ND0 U836 ( .I0(n1736), .I1(R[8]), .S(n512), .ZN(n515) );
  CKND2D0 U837 ( .A1(S[0]), .A2(n513), .ZN(n1039) );
  OAI222D0 U838 ( .A1(n1664), .A2(n1420), .B1(n1725), .B2(n1418), .C1(n1729), 
        .C2(n1728), .ZN(n517) );
  NR2D0 U839 ( .A1(n1736), .A2(n517), .ZN(n514) );
  CKND2D0 U840 ( .A1(n1039), .A2(n514), .ZN(n516) );
  AO21D0 U841 ( .A1(n515), .A2(n516), .B(\mult_x_9/n421 ), .Z(n1087) );
  CKND2D0 U842 ( .A1(R[8]), .A2(n517), .ZN(n518) );
  OAI221D0 U843 ( .A1(n518), .A2(n1039), .B1(R[8]), .B2(n517), .C(n516), .ZN(
        n1080) );
  INVD0 U844 ( .I(R[4]), .ZN(n596) );
  INVD0 U845 ( .I(R[3]), .ZN(n605) );
  AOI22D0 U846 ( .A1(R[3]), .A2(\mult_x_9/n686 ), .B1(R[2]), .B2(n605), .ZN(
        n525) );
  OAI22D0 U847 ( .A1(n596), .A2(n605), .B1(R[3]), .B2(R[4]), .ZN(n521) );
  ND3D0 U848 ( .A1(n519), .A2(n525), .A3(n521), .ZN(n1824) );
  INVD0 U849 ( .I(n525), .ZN(n520) );
  CKND2D0 U850 ( .A1(n520), .A2(n519), .ZN(n1740) );
  OAI22D0 U851 ( .A1(n1418), .A2(n1824), .B1(n1740), .B2(n1325), .ZN(n523) );
  OR2D0 U852 ( .A1(n519), .A2(n525), .Z(n1822) );
  OR2D0 U853 ( .A1(n521), .A2(n520), .Z(n1826) );
  OAI22D0 U854 ( .A1(n1726), .A2(n1822), .B1(n1728), .B2(n1826), .ZN(n522) );
  NR2D0 U855 ( .A1(n523), .A2(n522), .ZN(n524) );
  MUX2ND0 U856 ( .I0(\mult_x_9/n660 ), .I1(R[5]), .S(n524), .ZN(n1043) );
  NR2D0 U857 ( .A1(n1418), .A2(n525), .ZN(n1059) );
  NR2D0 U858 ( .A1(n1059), .A2(\mult_x_9/n660 ), .ZN(n526) );
  CKND2D0 U859 ( .A1(n526), .A2(n80), .ZN(n1042) );
  OR2D0 U860 ( .A1(n1043), .A2(n1042), .Z(n1040) );
  INVD0 U861 ( .I(n1740), .ZN(n1830) );
  NR2D0 U862 ( .A1(n1730), .A2(n1822), .ZN(n528) );
  OAI22D0 U863 ( .A1(n1726), .A2(n1826), .B1(n1728), .B2(n1824), .ZN(n527) );
  AOI211D0 U864 ( .A1(n1830), .A2(n1733), .B(n528), .C(n527), .ZN(n529) );
  MUX2ND0 U865 ( .I0(\mult_x_9/n660 ), .I1(R[5]), .S(n529), .ZN(n1041) );
  AO21D0 U866 ( .A1(n1039), .A2(n1040), .B(n1041), .Z(n1079) );
  AOI211D0 U867 ( .A1(n1723), .A2(n1830), .B(n531), .C(n530), .ZN(n532) );
  MUX2ND0 U868 ( .I0(\mult_x_9/n660 ), .I1(R[5]), .S(n532), .ZN(n1078) );
  NR2D0 U869 ( .A1(n1827), .A2(n1822), .ZN(n534) );
  AOI211D0 U870 ( .A1(n1719), .A2(n1830), .B(n534), .C(n533), .ZN(n535) );
  MUX2ND0 U871 ( .I0(\mult_x_9/n660 ), .I1(R[5]), .S(n535), .ZN(n1085) );
  INVD0 U872 ( .I(n536), .ZN(\mult_x_9/n419 ) );
  MUX2ND0 U873 ( .I0(R_lat_mag[11]), .I1(\mult_x_13/n608 ), .S(R_lat_mag[12]), 
        .ZN(n539) );
  NR2D0 U874 ( .A1(n1841), .A2(n539), .ZN(n1409) );
  MUX2ND0 U875 ( .I0(R_lat_mag[14]), .I1(n2028), .S(R_lat_mag[13]), .ZN(n540)
         );
  NR2D0 U876 ( .A1(n539), .A2(n540), .ZN(n2026) );
  INVD0 U877 ( .I(n2026), .ZN(n1962) );
  INVD0 U878 ( .I(R_lat_mag[12]), .ZN(n537) );
  MUX2ND0 U879 ( .I0(R_lat_mag[12]), .I1(n537), .S(R_lat_mag[13]), .ZN(n538)
         );
  IND2D0 U880 ( .A1(n538), .B1(n539), .ZN(n2021) );
  IND2D0 U881 ( .A1(n539), .B1(n540), .ZN(n2022) );
  OAI222D0 U882 ( .A1(n1962), .A2(n1843), .B1(n2021), .B2(n1841), .C1(n2174), 
        .C2(n2022), .ZN(n562) );
  OR3D0 U883 ( .A1(n1409), .A2(n2028), .A3(n562), .Z(n543) );
  IND3D0 U884 ( .A1(n540), .B1(n539), .B2(n538), .ZN(n2023) );
  OAI22D0 U885 ( .A1(n1841), .A2(n2023), .B1(n2170), .B2(n2022), .ZN(n541) );
  AOI211D0 U886 ( .A1(n2026), .A2(n1335), .B(n542), .C(n541), .ZN(n545) );
  CKND2D0 U887 ( .A1(R_lat_mag[14]), .A2(n545), .ZN(n544) );
  NR2D0 U888 ( .A1(n543), .A2(n544), .ZN(\mult_x_13/n388 ) );
  MUX2ND0 U889 ( .I0(R_lat_mag[8]), .I1(n2180), .S(R_lat_mag[9]), .ZN(n550) );
  NR2D0 U890 ( .A1(n1841), .A2(n550), .ZN(\mult_x_13/n418 ) );
  OAI211D0 U891 ( .A1(R_lat_mag[14]), .A2(n545), .B(n544), .C(n543), .ZN(n546)
         );
  IND2D0 U892 ( .A1(\mult_x_13/n388 ), .B1(n546), .ZN(n1370) );
  INVD0 U893 ( .I(R_lat_mag[9]), .ZN(n547) );
  MUX2ND0 U894 ( .I0(R_lat_mag[9]), .I1(n547), .S(R_lat_mag[10]), .ZN(n548) );
  MUX2ND0 U895 ( .I0(\mult_x_13/n608 ), .I1(R_lat_mag[11]), .S(R_lat_mag[10]), 
        .ZN(n551) );
  ND3D0 U896 ( .A1(n550), .A2(n548), .A3(n551), .ZN(n2032) );
  INVD0 U897 ( .I(n2032), .ZN(n2083) );
  INVD0 U898 ( .I(n550), .ZN(n549) );
  CKND2D0 U899 ( .A1(n549), .A2(n551), .ZN(n2030) );
  INVD0 U900 ( .I(n2030), .ZN(n2082) );
  AOI22D0 U901 ( .A1(inv_Q_mag[2]), .A2(n2083), .B1(n2167), .B2(n2082), .ZN(
        n553) );
  NR2D0 U902 ( .A1(n549), .A2(n548), .ZN(n2085) );
  NR2D0 U903 ( .A1(n551), .A2(n550), .ZN(n2084) );
  AOI22D0 U904 ( .A1(inv_Q_mag[3]), .A2(n2085), .B1(inv_Q_mag[4]), .B2(n2084), 
        .ZN(n552) );
  CKND2D0 U905 ( .A1(n553), .A2(n552), .ZN(n554) );
  MUX2ND0 U906 ( .I0(R_lat_mag[11]), .I1(\mult_x_13/n608 ), .S(n554), .ZN(
        n1362) );
  AOI22D0 U907 ( .A1(inv_Q_mag[0]), .A2(n2083), .B1(n1335), .B2(n2082), .ZN(
        n556) );
  AOI22D0 U908 ( .A1(inv_Q_mag[2]), .A2(n2084), .B1(inv_Q_mag[1]), .B2(n2085), 
        .ZN(n555) );
  CKND2D0 U909 ( .A1(n556), .A2(n555), .ZN(n1366) );
  NR2D0 U910 ( .A1(\mult_x_13/n608 ), .A2(n1366), .ZN(n1364) );
  AOI222D0 U911 ( .A1(n2082), .A2(n557), .B1(n2085), .B2(inv_Q_mag[0]), .C1(
        inv_Q_mag[1]), .C2(n2084), .ZN(n1838) );
  INVD0 U912 ( .I(n1838), .ZN(n1839) );
  NR3D0 U913 ( .A1(\mult_x_13/n418 ), .A2(\mult_x_13/n608 ), .A3(n1839), .ZN(
        n1365) );
  CKAN2D0 U914 ( .A1(n1364), .A2(n1365), .Z(n1408) );
  AOI22D0 U915 ( .A1(inv_Q_mag[1]), .A2(n2083), .B1(n2177), .B2(n2082), .ZN(
        n559) );
  AOI22D0 U916 ( .A1(inv_Q_mag[2]), .A2(n2085), .B1(inv_Q_mag[3]), .B2(n2084), 
        .ZN(n558) );
  CKND2D0 U917 ( .A1(n559), .A2(n558), .ZN(n560) );
  MUX2ND0 U918 ( .I0(\mult_x_13/n608 ), .I1(R_lat_mag[11]), .S(n560), .ZN(
        n1407) );
  OAI21D0 U919 ( .A1(n1408), .A2(n1409), .B(n1407), .ZN(n1361) );
  INVD0 U920 ( .I(n562), .ZN(n563) );
  CKND2D0 U921 ( .A1(R_lat_mag[14]), .A2(n1409), .ZN(n561) );
  MUX2ND0 U922 ( .I0(n563), .I1(n562), .S(n561), .ZN(n1360) );
  AOI22D0 U923 ( .A1(inv_Q_mag[3]), .A2(n2083), .B1(n2162), .B2(n2082), .ZN(
        n565) );
  CKND2D0 U924 ( .A1(n565), .A2(n564), .ZN(n566) );
  MUX2ND0 U925 ( .I0(R_lat_mag[11]), .I1(\mult_x_13/n608 ), .S(n566), .ZN(
        n1368) );
  INVD0 U926 ( .I(n567), .ZN(\mult_x_13/n386 ) );
  FA1D0 U927 ( .A(n570), .B(n569), .CI(n568), .CO(n571), .S(n167) );
  INVD0 U928 ( .I(n571), .ZN(\mult_x_13/n419 ) );
  OAI22D0 U929 ( .A1(n768), .A2(n1477), .B1(R[20]), .B2(R[21]), .ZN(n1379) );
  NR2D0 U930 ( .A1(n1379), .A2(R[22]), .ZN(n1322) );
  INVD0 U931 ( .I(n1322), .ZN(n1417) );
  INVD0 U932 ( .I(S[19]), .ZN(n1757) );
  INVD0 U933 ( .I(R[22]), .ZN(n800) );
  AOI33D0 U934 ( .A1(R[22]), .A2(n768), .A3(n1477), .B1(R[21]), .B2(R[20]), 
        .B3(n800), .ZN(n1419) );
  INVD0 U935 ( .I(n1419), .ZN(n1384) );
  ND3D0 U936 ( .A1(R[22]), .A2(R[21]), .A3(R[20]), .ZN(n1394) );
  INVD0 U937 ( .I(n1394), .ZN(n1383) );
  AOI22D0 U938 ( .A1(S[18]), .A2(n1384), .B1(S[17]), .B2(n1383), .ZN(n574) );
  FA1D0 U939 ( .A(S[4]), .B(S[5]), .CI(n572), .CO(n988), .S(n1719) );
  NR2D0 U940 ( .A1(n800), .A2(n1379), .ZN(n1385) );
  CKND2D0 U941 ( .A1(n1760), .A2(n1385), .ZN(n573) );
  OAI211D0 U942 ( .A1(n1417), .A2(n1757), .B(n574), .C(n573), .ZN(
        \mult_x_9/n511 ) );
  INVD0 U943 ( .I(S[13]), .ZN(n1787) );
  AOI22D0 U944 ( .A1(S[12]), .A2(n1384), .B1(S[11]), .B2(n1383), .ZN(n577) );
  FA1D0 U945 ( .A(S[12]), .B(S[13]), .CI(n575), .CO(n940), .S(n1790) );
  CKND2D0 U946 ( .A1(n1790), .A2(n1385), .ZN(n576) );
  OAI211D0 U947 ( .A1(n1417), .A2(n1787), .B(n577), .C(n576), .ZN(
        \mult_x_9/n517 ) );
  AOI22D0 U948 ( .A1(S[6]), .A2(n1384), .B1(S[5]), .B2(n1383), .ZN(n580) );
  FA1D0 U949 ( .A(S[6]), .B(S[7]), .CI(n578), .CO(n1011), .S(n1820) );
  CKND2D0 U950 ( .A1(n1820), .A2(n1385), .ZN(n579) );
  OAI211D0 U951 ( .A1(n1417), .A2(n1817), .B(n580), .C(n579), .ZN(
        \mult_x_9/n522 ) );
  INVD0 U952 ( .I(inv_Q_mag[13]), .ZN(n2127) );
  INVD0 U953 ( .I(n1842), .ZN(n1336) );
  AOI22D0 U954 ( .A1(inv_Q_mag[12]), .A2(n1336), .B1(n2226), .B2(n1334), .ZN(
        n582) );
  CKND2D0 U955 ( .A1(inv_Q_mag[11]), .A2(n1337), .ZN(n581) );
  OAI211D0 U956 ( .A1(n1840), .A2(n2127), .B(n582), .C(n581), .ZN(
        \mult_x_13/n517 ) );
  AOI22D0 U957 ( .A1(inv_Q_mag[6]), .A2(n1336), .B1(n2250), .B2(n1334), .ZN(
        n584) );
  CKND2D0 U958 ( .A1(inv_Q_mag[5]), .A2(n1337), .ZN(n583) );
  OAI211D0 U959 ( .A1(n1840), .A2(n2151), .B(n584), .C(n583), .ZN(
        \mult_x_13/n522 ) );
  AOI22D0 U960 ( .A1(inv_Q_mag[18]), .A2(n1336), .B1(inv_Q_mag[17]), .B2(n1337), .ZN(n586) );
  CKND2D0 U961 ( .A1(n2202), .A2(n1334), .ZN(n585) );
  OAI211D0 U962 ( .A1(n1840), .A2(n2103), .B(n586), .C(n585), .ZN(
        \mult_x_13/n511 ) );
  IND2D0 U963 ( .A1(n601), .B1(n1726), .ZN(n1053) );
  OR2D0 U964 ( .A1(n1053), .A2(S[3]), .Z(n606) );
  CKND2D0 U965 ( .A1(n592), .A2(n1827), .ZN(n590) );
  NR2D0 U966 ( .A1(S[6]), .A2(n590), .ZN(n613) );
  INVD0 U967 ( .I(S[23]), .ZN(n1388) );
  OR2D0 U968 ( .A1(n613), .A2(n1388), .Z(n587) );
  MUX2ND0 U969 ( .I0(S[7]), .I1(n1817), .S(n587), .ZN(n618) );
  CKND2D0 U970 ( .A1(n1047), .A2(\mult_x_9/n686 ), .ZN(n603) );
  NR2D0 U971 ( .A1(R[3]), .A2(n603), .ZN(n594) );
  CKND2D0 U972 ( .A1(n594), .A2(n596), .ZN(n608) );
  IND2D0 U973 ( .A1(n608), .B1(\mult_x_9/n660 ), .ZN(n610) );
  CKND2D0 U974 ( .A1(R[23]), .A2(n610), .ZN(n588) );
  MUX2ND0 U975 ( .I0(R[6]), .I1(n589), .S(n588), .ZN(n654) );
  INVD0 U976 ( .I(S[6]), .ZN(n1823) );
  CKND2D0 U977 ( .A1(S[23]), .A2(n590), .ZN(n591) );
  MUX2ND0 U978 ( .I0(n1823), .I1(S[6]), .S(n591), .ZN(n621) );
  OR2D0 U979 ( .A1(n592), .A2(n1388), .Z(n593) );
  MUX2ND0 U980 ( .I0(S[5]), .I1(n1827), .S(n593), .ZN(n624) );
  INVD0 U981 ( .I(R[23]), .ZN(n1389) );
  NR2D0 U982 ( .A1(n594), .A2(n1389), .ZN(n595) );
  MUX2ND0 U983 ( .I0(n596), .I1(R[4]), .S(n595), .ZN(n650) );
  CKND2D0 U984 ( .A1(S[23]), .A2(n1053), .ZN(n597) );
  MUX2ND0 U985 ( .I0(S[3]), .I1(n1730), .S(n597), .ZN(n630) );
  NR2D0 U986 ( .A1(n1047), .A2(n1389), .ZN(n598) );
  MUX2ND0 U987 ( .I0(\mult_x_9/n686 ), .I1(R[2]), .S(n598), .ZN(n646) );
  NR2D0 U988 ( .A1(R[0]), .A2(n1418), .ZN(n636) );
  OAI32D0 U989 ( .A1(n1388), .A2(n1728), .A3(n1418), .B1(S[1]), .B2(S[23]), 
        .ZN(n643) );
  INVD0 U990 ( .I(n643), .ZN(n600) );
  CKND2D0 U991 ( .A1(n601), .A2(n600), .ZN(n644) );
  INVD0 U992 ( .I(n644), .ZN(n637) );
  INVD0 U993 ( .I(R[1]), .ZN(n1044) );
  CKND2D0 U994 ( .A1(R[23]), .A2(R[0]), .ZN(n599) );
  MUX2ND0 U995 ( .I0(n1044), .I1(R[1]), .S(n599), .ZN(n645) );
  OAI222D0 U996 ( .A1(n636), .A2(n637), .B1(n636), .B2(n645), .C1(n645), .C2(
        n600), .ZN(n635) );
  CKND2D0 U997 ( .A1(S[23]), .A2(n601), .ZN(n602) );
  MUX2ND0 U998 ( .I0(n1726), .I1(S[2]), .S(n602), .ZN(n633) );
  MAOI222D0 U999 ( .A(n646), .B(n635), .C(n633), .ZN(n632) );
  CKND2D0 U1000 ( .A1(R[23]), .A2(n603), .ZN(n604) );
  MUX2ND0 U1001 ( .I0(n605), .I1(R[3]), .S(n604), .ZN(n649) );
  MAOI222D0 U1002 ( .A(n630), .B(n632), .C(n649), .ZN(n628) );
  CKND2D0 U1003 ( .A1(S[23]), .A2(n606), .ZN(n607) );
  MUX2ND0 U1004 ( .I0(n1825), .I1(S[4]), .S(n607), .ZN(n627) );
  MAOI222D0 U1005 ( .A(n650), .B(n628), .C(n627), .ZN(n626) );
  CKND2D0 U1006 ( .A1(R[23]), .A2(n608), .ZN(n609) );
  MUX2ND0 U1007 ( .I0(\mult_x_9/n660 ), .I1(R[5]), .S(n609), .ZN(n652) );
  MAOI222D0 U1008 ( .A(n624), .B(n626), .C(n652), .ZN(n622) );
  MAOI222D0 U1009 ( .A(n654), .B(n621), .C(n622), .ZN(n620) );
  NR2D0 U1010 ( .A1(n610), .A2(R[6]), .ZN(n615) );
  NR2D0 U1011 ( .A1(n615), .A2(n1389), .ZN(n611) );
  MUX2ND0 U1012 ( .I0(R[7]), .I1(n612), .S(n611), .ZN(n656) );
  MAOI222D0 U1013 ( .A(n618), .B(n620), .C(n656), .ZN(n703) );
  INVD0 U1014 ( .I(n703), .ZN(n617) );
  INVD0 U1015 ( .I(S[8]), .ZN(n1812) );
  CKND2D0 U1016 ( .A1(n613), .A2(n1817), .ZN(n659) );
  CKND2D0 U1017 ( .A1(S[23]), .A2(n659), .ZN(n614) );
  MUX2ND0 U1018 ( .I0(n1812), .I1(S[8]), .S(n614), .ZN(n704) );
  INVD0 U1019 ( .I(n704), .ZN(n658) );
  INR2D0 U1020 ( .A1(n615), .B1(R[7]), .ZN(n661) );
  NR2D0 U1021 ( .A1(n661), .A2(n1389), .ZN(n616) );
  MUX2ND0 U1022 ( .I0(n1736), .I1(R[8]), .S(n616), .ZN(n705) );
  MUX2ND0 U1023 ( .I0(n658), .I1(n704), .S(n705), .ZN(n665) );
  MUX2ND0 U1024 ( .I0(n617), .I1(n703), .S(n665), .ZN(sub_tc[8]) );
  INVD0 U1025 ( .I(n620), .ZN(n619) );
  INVD0 U1026 ( .I(n618), .ZN(n657) );
  MUX2ND0 U1027 ( .I0(n657), .I1(n618), .S(n656), .ZN(n685) );
  MUX2ND0 U1028 ( .I0(n620), .I1(n619), .S(n685), .ZN(sub_tc[7]) );
  INVD0 U1029 ( .I(n622), .ZN(n623) );
  INVD0 U1030 ( .I(n621), .ZN(n655) );
  MUX2ND0 U1031 ( .I0(n655), .I1(n621), .S(n654), .ZN(n668) );
  MUX2ND0 U1032 ( .I0(n623), .I1(n622), .S(n668), .ZN(sub_tc[6]) );
  INVD0 U1033 ( .I(n626), .ZN(n625) );
  INVD0 U1034 ( .I(n624), .ZN(n653) );
  MUX2ND0 U1035 ( .I0(n653), .I1(n624), .S(n652), .ZN(n682) );
  MUX2ND0 U1036 ( .I0(n626), .I1(n625), .S(n682), .ZN(sub_tc[5]) );
  INVD0 U1037 ( .I(n628), .ZN(n629) );
  INVD0 U1038 ( .I(n627), .ZN(n651) );
  MUX2ND0 U1039 ( .I0(n651), .I1(n627), .S(n650), .ZN(n671) );
  MUX2ND0 U1040 ( .I0(n629), .I1(n628), .S(n671), .ZN(sub_tc[4]) );
  INVD0 U1041 ( .I(n632), .ZN(n631) );
  INVD0 U1042 ( .I(n630), .ZN(n648) );
  MUX2ND0 U1043 ( .I0(n648), .I1(n630), .S(n649), .ZN(n674) );
  MUX2ND0 U1044 ( .I0(n632), .I1(n631), .S(n674), .ZN(sub_tc[3]) );
  INVD0 U1045 ( .I(n635), .ZN(n634) );
  INVD0 U1046 ( .I(n633), .ZN(n647) );
  MUX2ND0 U1047 ( .I0(n633), .I1(n647), .S(n646), .ZN(n677) );
  MUX2ND0 U1048 ( .I0(n635), .I1(n634), .S(n677), .ZN(sub_tc[2]) );
  INVD0 U1049 ( .I(n636), .ZN(n641) );
  INVD0 U1050 ( .I(sub_tc[7]), .ZN(n639) );
  INVD0 U1051 ( .I(sub_tc[5]), .ZN(n906) );
  INVD0 U1052 ( .I(sub_tc[3]), .ZN(n929) );
  INVD0 U1053 ( .I(add_tc[0]), .ZN(n921) );
  MUX2ND0 U1054 ( .I0(n637), .I1(n644), .S(n645), .ZN(n681) );
  CKND2D0 U1055 ( .A1(n681), .A2(n641), .ZN(n640) );
  CKND2D0 U1056 ( .A1(n921), .A2(n640), .ZN(n807) );
  NR2D0 U1057 ( .A1(sub_tc[2]), .A2(n807), .ZN(n928) );
  CKND2D0 U1058 ( .A1(n929), .A2(n928), .ZN(n927) );
  NR2D0 U1059 ( .A1(sub_tc[4]), .A2(n927), .ZN(n912) );
  CKND2D0 U1060 ( .A1(n906), .A2(n912), .ZN(n905) );
  NR2D0 U1061 ( .A1(sub_tc[6]), .A2(n905), .ZN(n867) );
  CKND2D0 U1062 ( .A1(n639), .A2(n867), .ZN(n638) );
  AOI21D0 U1063 ( .A1(sub_tc[8]), .A2(n638), .B(n870), .ZN(N133) );
  OAI21D0 U1064 ( .A1(n681), .A2(n641), .B(n640), .ZN(sub_tc[1]) );
  CKND2D0 U1065 ( .A1(R[0]), .A2(S[0]), .ZN(n680) );
  OAI222D0 U1066 ( .A1(n645), .A2(n644), .B1(n645), .B2(n680), .C1(n680), .C2(
        n643), .ZN(n678) );
  MAOI222D0 U1067 ( .A(n647), .B(n646), .C(n678), .ZN(n675) );
  MAOI222D0 U1068 ( .A(n649), .B(n648), .C(n675), .ZN(n673) );
  MAOI222D0 U1069 ( .A(n651), .B(n650), .C(n673), .ZN(n683) );
  MAOI222D0 U1070 ( .A(n683), .B(n653), .C(n652), .ZN(n670) );
  MAOI222D0 U1071 ( .A(n655), .B(n654), .C(n670), .ZN(n686) );
  MAOI222D0 U1072 ( .A(n686), .B(n657), .C(n656), .ZN(n667) );
  MAOI222D0 U1073 ( .A(n658), .B(n705), .C(n667), .ZN(n810) );
  INVD0 U1074 ( .I(n810), .ZN(n664) );
  INVD0 U1075 ( .I(S[9]), .ZN(n1807) );
  NR2D0 U1076 ( .A1(S[8]), .A2(n659), .ZN(n689) );
  OR2D0 U1077 ( .A1(n689), .A2(n1388), .Z(n660) );
  MUX2ND0 U1078 ( .I0(S[9]), .I1(n1807), .S(n660), .ZN(n706) );
  INVD0 U1079 ( .I(n706), .ZN(n809) );
  CKND2D0 U1080 ( .A1(R[23]), .A2(n691), .ZN(n662) );
  MUX2ND0 U1081 ( .I0(n663), .I1(R[9]), .S(n662), .ZN(n808) );
  MUX2ND0 U1082 ( .I0(n706), .I1(n809), .S(n808), .ZN(n723) );
  MUX2ND0 U1083 ( .I0(n810), .I1(n664), .S(n723), .ZN(add_tc[9]) );
  INVD0 U1084 ( .I(n667), .ZN(n666) );
  MUX2ND0 U1085 ( .I0(n667), .I1(n666), .S(n665), .ZN(add_tc[8]) );
  INVD0 U1086 ( .I(n670), .ZN(n669) );
  MUX2ND0 U1087 ( .I0(n670), .I1(n669), .S(n668), .ZN(add_tc[6]) );
  INVD0 U1088 ( .I(n673), .ZN(n672) );
  MUX2ND0 U1089 ( .I0(n673), .I1(n672), .S(n671), .ZN(add_tc[4]) );
  INVD0 U1090 ( .I(n675), .ZN(n676) );
  MUX2ND0 U1091 ( .I0(n676), .I1(n675), .S(n674), .ZN(add_tc[3]) );
  MUX2ND0 U1092 ( .I0(n679), .I1(n678), .S(n677), .ZN(add_tc[2]) );
  CKND2D0 U1093 ( .A1(n681), .A2(n680), .ZN(n920) );
  OAI21D0 U1094 ( .A1(n681), .A2(n680), .B(n920), .ZN(add_tc[1]) );
  INVD0 U1095 ( .I(n683), .ZN(n684) );
  MUX2ND0 U1096 ( .I0(n684), .I1(n683), .S(n682), .ZN(add_tc[5]) );
  INVD0 U1097 ( .I(n686), .ZN(n687) );
  MUX2ND0 U1098 ( .I0(n687), .I1(n686), .S(n685), .ZN(add_tc[7]) );
  INVD0 U1099 ( .I(add_tc[9]), .ZN(n688) );
  INVD0 U1100 ( .I(add_tc[3]), .ZN(n911) );
  OR2D0 U1101 ( .A1(add_tc[1]), .A2(add_tc[0]), .Z(n919) );
  NR2D0 U1102 ( .A1(add_tc[2]), .A2(n919), .ZN(n913) );
  NR2D0 U1103 ( .A1(add_tc[4]), .A2(n923), .ZN(n922) );
  INVD0 U1104 ( .I(add_tc[5]), .ZN(n902) );
  CKND2D0 U1105 ( .A1(n922), .A2(n902), .ZN(n901) );
  NR2D0 U1106 ( .A1(add_tc[6]), .A2(n901), .ZN(n909) );
  INVD0 U1107 ( .I(add_tc[7]), .ZN(n908) );
  CKND2D0 U1108 ( .A1(n909), .A2(n908), .ZN(n907) );
  NR2D0 U1109 ( .A1(add_tc[8]), .A2(n907), .ZN(n804) );
  CKND2D0 U1110 ( .A1(n688), .A2(n804), .ZN(n878) );
  OA21D0 U1111 ( .A1(n688), .A2(n804), .B(n878), .Z(N83) );
  CKND2D0 U1112 ( .A1(n689), .A2(n1807), .ZN(n701) );
  NR2D0 U1113 ( .A1(S[10]), .A2(n701), .ZN(n696) );
  INVD0 U1114 ( .I(S[11]), .ZN(n1797) );
  CKND2D0 U1115 ( .A1(n696), .A2(n1797), .ZN(n694) );
  NR2D0 U1116 ( .A1(S[12]), .A2(n694), .ZN(n712) );
  OR2D0 U1117 ( .A1(n712), .A2(n1388), .Z(n690) );
  MUX2ND0 U1118 ( .I0(S[13]), .I1(n1787), .S(n690), .ZN(n729) );
  NR2D0 U1119 ( .A1(R[9]), .A2(n691), .ZN(n698) );
  CKND2D0 U1120 ( .A1(\mult_x_9/n608 ), .A2(n707), .ZN(n709) );
  CKND2D0 U1121 ( .A1(R[23]), .A2(n709), .ZN(n692) );
  MUX2ND0 U1122 ( .I0(R[12]), .I1(n693), .S(n692), .ZN(n815) );
  INVD0 U1123 ( .I(S[12]), .ZN(n1792) );
  CKND2D0 U1124 ( .A1(S[23]), .A2(n694), .ZN(n695) );
  MUX2ND0 U1125 ( .I0(n1792), .I1(S[12]), .S(n695), .ZN(n717) );
  OR2D0 U1126 ( .A1(n696), .A2(n1388), .Z(n697) );
  MUX2ND0 U1127 ( .I0(S[11]), .I1(n1797), .S(n697), .ZN(n726) );
  NR2D0 U1128 ( .A1(n698), .A2(n1389), .ZN(n699) );
  MUX2ND0 U1129 ( .I0(n700), .I1(R[10]), .S(n699), .ZN(n811) );
  INVD0 U1130 ( .I(S[10]), .ZN(n1802) );
  CKND2D0 U1131 ( .A1(S[23]), .A2(n701), .ZN(n702) );
  MUX2ND0 U1132 ( .I0(n1802), .I1(S[10]), .S(n702), .ZN(n720) );
  MAOI222D0 U1133 ( .A(n705), .B(n704), .C(n703), .ZN(n724) );
  MAOI222D0 U1134 ( .A(n706), .B(n724), .C(n808), .ZN(n722) );
  MAOI222D0 U1135 ( .A(n811), .B(n720), .C(n722), .ZN(n727) );
  NR2D0 U1136 ( .A1(n707), .A2(n1389), .ZN(n708) );
  MUX2ND0 U1137 ( .I0(R[11]), .I1(\mult_x_9/n608 ), .S(n708), .ZN(n813) );
  MAOI222D0 U1138 ( .A(n726), .B(n727), .C(n813), .ZN(n719) );
  MAOI222D0 U1139 ( .A(n815), .B(n717), .C(n719), .ZN(n730) );
  NR2D0 U1140 ( .A1(n709), .A2(R[12]), .ZN(n714) );
  MUX2ND0 U1141 ( .I0(R[13]), .I1(n711), .S(n710), .ZN(n817) );
  MAOI222D0 U1142 ( .A(n729), .B(n730), .C(n817), .ZN(n756) );
  INVD0 U1143 ( .I(S[14]), .ZN(n1782) );
  CKND2D0 U1144 ( .A1(S[23]), .A2(n734), .ZN(n713) );
  MUX2ND0 U1145 ( .I0(n1782), .I1(S[14]), .S(n713), .ZN(n757) );
  INVD0 U1146 ( .I(n757), .ZN(n820) );
  INR2D0 U1147 ( .A1(n714), .B1(R[13]), .ZN(n736) );
  NR2D0 U1148 ( .A1(n736), .A2(n1389), .ZN(n715) );
  MUX2ND0 U1149 ( .I0(n1603), .I1(R[14]), .S(n715), .ZN(n819) );
  MUX2ND0 U1150 ( .I0(n757), .I1(n820), .S(n819), .ZN(n852) );
  MUX2ND0 U1151 ( .I0(n756), .I1(n716), .S(n852), .ZN(sub_tc[14]) );
  INVD0 U1152 ( .I(n719), .ZN(n718) );
  INVD0 U1153 ( .I(n717), .ZN(n816) );
  MUX2ND0 U1154 ( .I0(n717), .I1(n816), .S(n815), .ZN(n858) );
  MUX2ND0 U1155 ( .I0(n719), .I1(n718), .S(n858), .ZN(sub_tc[12]) );
  INVD0 U1156 ( .I(n722), .ZN(n721) );
  INVD0 U1157 ( .I(n720), .ZN(n812) );
  MUX2ND0 U1158 ( .I0(n720), .I1(n812), .S(n811), .ZN(n864) );
  MUX2ND0 U1159 ( .I0(n722), .I1(n721), .S(n864), .ZN(sub_tc[10]) );
  INVD0 U1160 ( .I(n724), .ZN(n725) );
  MUX2ND0 U1161 ( .I0(n725), .I1(n724), .S(n723), .ZN(sub_tc[9]) );
  INVD0 U1162 ( .I(n727), .ZN(n728) );
  INVD0 U1163 ( .I(n726), .ZN(n814) );
  MUX2ND0 U1164 ( .I0(n726), .I1(n814), .S(n813), .ZN(n861) );
  MUX2ND0 U1165 ( .I0(n728), .I1(n727), .S(n861), .ZN(sub_tc[11]) );
  INVD0 U1166 ( .I(n730), .ZN(n731) );
  INVD0 U1167 ( .I(n729), .ZN(n818) );
  MUX2ND0 U1168 ( .I0(n729), .I1(n818), .S(n817), .ZN(n855) );
  MUX2ND0 U1169 ( .I0(n731), .I1(n730), .S(n855), .ZN(sub_tc[13]) );
  INVD0 U1170 ( .I(sub_tc[9]), .ZN(n869) );
  CKND2D0 U1171 ( .A1(n870), .A2(n869), .ZN(n900) );
  NR2D0 U1172 ( .A1(sub_tc[10]), .A2(n900), .ZN(n899) );
  INVD0 U1173 ( .I(sub_tc[11]), .ZN(n797) );
  CKND2D0 U1174 ( .A1(n899), .A2(n797), .ZN(n796) );
  NR2D0 U1175 ( .A1(sub_tc[12]), .A2(n796), .ZN(n795) );
  INVD0 U1176 ( .I(sub_tc[13]), .ZN(n733) );
  CKND2D0 U1177 ( .A1(n795), .A2(n733), .ZN(n732) );
  NR2D0 U1178 ( .A1(sub_tc[14]), .A2(n732), .ZN(n806) );
  AOI21D0 U1179 ( .A1(sub_tc[14]), .A2(n732), .B(n806), .ZN(N139) );
  OA21D0 U1180 ( .A1(n795), .A2(n733), .B(n732), .Z(N138) );
  INVD0 U1181 ( .I(S[21]), .ZN(n1747) );
  NR2D0 U1182 ( .A1(S[14]), .A2(n734), .ZN(n754) );
  INVD0 U1183 ( .I(S[15]), .ZN(n1777) );
  CKND2D0 U1184 ( .A1(n754), .A2(n1777), .ZN(n752) );
  NR2D0 U1185 ( .A1(S[16]), .A2(n752), .ZN(n747) );
  INVD0 U1186 ( .I(S[17]), .ZN(n1767) );
  CKND2D0 U1187 ( .A1(n747), .A2(n1767), .ZN(n745) );
  NR2D0 U1188 ( .A1(S[18]), .A2(n745), .ZN(n740) );
  CKND2D0 U1189 ( .A1(n740), .A2(n1757), .ZN(n738) );
  NR2D0 U1190 ( .A1(S[20]), .A2(n738), .ZN(n769) );
  OR2D0 U1191 ( .A1(n769), .A2(n1388), .Z(n735) );
  MUX2ND0 U1192 ( .I0(S[21]), .I1(n1747), .S(n735), .ZN(n792) );
  CKND2D0 U1193 ( .A1(n736), .A2(n1603), .ZN(n758) );
  NR2D0 U1194 ( .A1(R[15]), .A2(n758), .ZN(n749) );
  CKND2D0 U1195 ( .A1(\mult_x_9/n556 ), .A2(n761), .ZN(n742) );
  NR2D0 U1196 ( .A1(n742), .A2(R[18]), .ZN(n763) );
  INR2D0 U1197 ( .A1(n763), .B1(R[19]), .ZN(n766) );
  NR2D0 U1198 ( .A1(n766), .A2(n1389), .ZN(n737) );
  MUX2ND0 U1199 ( .I0(n1477), .I1(R[20]), .S(n737), .ZN(n831) );
  INVD0 U1200 ( .I(S[20]), .ZN(n1752) );
  CKND2D0 U1201 ( .A1(S[23]), .A2(n738), .ZN(n739) );
  MUX2ND0 U1202 ( .I0(n1752), .I1(S[20]), .S(n739), .ZN(n774) );
  OR2D0 U1203 ( .A1(n740), .A2(n1388), .Z(n741) );
  MUX2ND0 U1204 ( .I0(S[19]), .I1(n1757), .S(n741), .ZN(n789) );
  CKND2D0 U1205 ( .A1(R[23]), .A2(n742), .ZN(n743) );
  MUX2ND0 U1206 ( .I0(R[18]), .I1(n744), .S(n743), .ZN(n827) );
  INVD0 U1207 ( .I(S[18]), .ZN(n1762) );
  CKND2D0 U1208 ( .A1(S[23]), .A2(n745), .ZN(n746) );
  MUX2ND0 U1209 ( .I0(n1762), .I1(S[18]), .S(n746), .ZN(n777) );
  OR2D0 U1210 ( .A1(n747), .A2(n1388), .Z(n748) );
  MUX2ND0 U1211 ( .I0(S[17]), .I1(n1767), .S(n748), .ZN(n786) );
  NR2D0 U1212 ( .A1(n749), .A2(n1389), .ZN(n750) );
  MUX2ND0 U1213 ( .I0(n751), .I1(R[16]), .S(n750), .ZN(n823) );
  INVD0 U1214 ( .I(S[16]), .ZN(n1772) );
  MUX2ND0 U1215 ( .I0(n1772), .I1(S[16]), .S(n753), .ZN(n780) );
  OR2D0 U1216 ( .A1(n754), .A2(n1388), .Z(n755) );
  MUX2ND0 U1217 ( .I0(S[15]), .I1(n1777), .S(n755), .ZN(n783) );
  MAOI222D0 U1218 ( .A(n819), .B(n757), .C(n756), .ZN(n784) );
  CKND2D0 U1219 ( .A1(R[23]), .A2(n758), .ZN(n759) );
  MUX2ND0 U1220 ( .I0(n760), .I1(R[15]), .S(n759), .ZN(n821) );
  MAOI222D0 U1221 ( .A(n783), .B(n784), .C(n821), .ZN(n782) );
  MAOI222D0 U1222 ( .A(n823), .B(n780), .C(n782), .ZN(n787) );
  NR2D0 U1223 ( .A1(n761), .A2(n1389), .ZN(n762) );
  MUX2ND0 U1224 ( .I0(R[17]), .I1(\mult_x_9/n556 ), .S(n762), .ZN(n825) );
  MAOI222D0 U1225 ( .A(n786), .B(n787), .C(n825), .ZN(n779) );
  MAOI222D0 U1226 ( .A(n827), .B(n777), .C(n779), .ZN(n790) );
  MUX2ND0 U1227 ( .I0(R[19]), .I1(n765), .S(n764), .ZN(n829) );
  MAOI222D0 U1228 ( .A(n789), .B(n790), .C(n829), .ZN(n776) );
  MAOI222D0 U1229 ( .A(n831), .B(n774), .C(n776), .ZN(n793) );
  CKND2D0 U1230 ( .A1(R[23]), .A2(n771), .ZN(n767) );
  MUX2ND0 U1231 ( .I0(n768), .I1(R[21]), .S(n767), .ZN(n833) );
  MAOI222D0 U1232 ( .A(n792), .B(n793), .C(n833), .ZN(n799) );
  INVD0 U1233 ( .I(S[22]), .ZN(n1742) );
  CKND2D0 U1234 ( .A1(n769), .A2(n1747), .ZN(n802) );
  CKND2D0 U1235 ( .A1(S[23]), .A2(n802), .ZN(n770) );
  MUX2ND0 U1236 ( .I0(n1742), .I1(S[22]), .S(n770), .ZN(n798) );
  NR2D0 U1237 ( .A1(R[21]), .A2(n771), .ZN(n801) );
  NR2D0 U1238 ( .A1(n801), .A2(n1389), .ZN(n772) );
  MUX2ND0 U1239 ( .I0(n800), .I1(R[22]), .S(n772), .ZN(n835) );
  MUX2ND0 U1240 ( .I0(n798), .I1(n836), .S(n835), .ZN(n884) );
  MUX2ND0 U1241 ( .I0(n799), .I1(n773), .S(n884), .ZN(sub_tc[22]) );
  INVD0 U1242 ( .I(n776), .ZN(n775) );
  INVD0 U1243 ( .I(n774), .ZN(n832) );
  MUX2ND0 U1244 ( .I0(n774), .I1(n832), .S(n831), .ZN(n871) );
  MUX2ND0 U1245 ( .I0(n776), .I1(n775), .S(n871), .ZN(sub_tc[20]) );
  INVD0 U1246 ( .I(n779), .ZN(n778) );
  INVD0 U1247 ( .I(n777), .ZN(n828) );
  MUX2ND0 U1248 ( .I0(n777), .I1(n828), .S(n827), .ZN(n840) );
  MUX2ND0 U1249 ( .I0(n779), .I1(n778), .S(n840), .ZN(sub_tc[18]) );
  INVD0 U1250 ( .I(n782), .ZN(n781) );
  INVD0 U1251 ( .I(n780), .ZN(n824) );
  MUX2ND0 U1252 ( .I0(n780), .I1(n824), .S(n823), .ZN(n846) );
  MUX2ND0 U1253 ( .I0(n782), .I1(n781), .S(n846), .ZN(sub_tc[16]) );
  INVD0 U1254 ( .I(n784), .ZN(n785) );
  INVD0 U1255 ( .I(n783), .ZN(n822) );
  MUX2ND0 U1256 ( .I0(n783), .I1(n822), .S(n821), .ZN(n849) );
  MUX2ND0 U1257 ( .I0(n785), .I1(n784), .S(n849), .ZN(sub_tc[15]) );
  INVD0 U1258 ( .I(n786), .ZN(n826) );
  MUX2ND0 U1259 ( .I0(n786), .I1(n826), .S(n825), .ZN(n843) );
  MUX2ND0 U1260 ( .I0(n788), .I1(n787), .S(n843), .ZN(sub_tc[17]) );
  INVD0 U1261 ( .I(n790), .ZN(n791) );
  INVD0 U1262 ( .I(n789), .ZN(n830) );
  MUX2ND0 U1263 ( .I0(n789), .I1(n830), .S(n829), .ZN(n874) );
  MUX2ND0 U1264 ( .I0(n791), .I1(n790), .S(n874), .ZN(sub_tc[19]) );
  INVD0 U1265 ( .I(n793), .ZN(n794) );
  INVD0 U1266 ( .I(n792), .ZN(n834) );
  MUX2ND0 U1267 ( .I0(n792), .I1(n834), .S(n833), .ZN(n887) );
  MUX2ND0 U1268 ( .I0(n794), .I1(n793), .S(n887), .ZN(sub_tc[21]) );
  INVD0 U1269 ( .I(sub_tc[15]), .ZN(n805) );
  CKND2D0 U1270 ( .A1(n806), .A2(n805), .ZN(n883) );
  NR2D0 U1271 ( .A1(sub_tc[16]), .A2(n883), .ZN(n882) );
  INVD0 U1272 ( .I(sub_tc[17]), .ZN(n839) );
  CKND2D0 U1273 ( .A1(n882), .A2(n839), .ZN(n918) );
  INVD0 U1274 ( .I(sub_tc[19]), .ZN(n904) );
  CKND2D0 U1275 ( .A1(n917), .A2(n904), .ZN(n903) );
  NR2D0 U1276 ( .A1(sub_tc[20]), .A2(n903), .ZN(n895) );
  INVD0 U1277 ( .I(sub_tc[21]), .ZN(n894) );
  CKND2D0 U1278 ( .A1(n895), .A2(n894), .ZN(n893) );
  NR2D0 U1279 ( .A1(sub_tc[22]), .A2(n893), .ZN(n2264) );
  AOI21D0 U1280 ( .A1(sub_tc[22]), .A2(n893), .B(n2264), .ZN(N147) );
  AOI21D0 U1281 ( .A1(sub_tc[12]), .A2(n796), .B(n795), .ZN(N137) );
  OA21D0 U1282 ( .A1(n899), .A2(n797), .B(n796), .Z(N136) );
  MAOI222D0 U1283 ( .A(n835), .B(n799), .C(n798), .ZN(n803) );
  AOI21D0 U1284 ( .A1(n801), .A2(n800), .B(n1389), .ZN(n933) );
  INVD0 U1285 ( .I(n933), .ZN(n931) );
  OAI21D0 U1286 ( .A1(S[22]), .A2(n802), .B(S[23]), .ZN(n932) );
  CKXOR2D0 U1287 ( .A1(n931), .A2(n932), .Z(n837) );
  NR2D0 U1288 ( .A1(n803), .A2(n837), .ZN(n934) );
  AOI21D0 U1289 ( .A1(n803), .A2(n837), .B(n934), .ZN(sub_tc[23]) );
  AOI21D0 U1290 ( .A1(add_tc[8]), .A2(n907), .B(n804), .ZN(N82) );
  OA21D0 U1291 ( .A1(n806), .A2(n805), .B(n883), .Z(N140) );
  AOI21D0 U1292 ( .A1(sub_tc[2]), .A2(n807), .B(n928), .ZN(N127) );
  MAOI222D0 U1293 ( .A(n810), .B(n809), .C(n808), .ZN(n865) );
  MAOI222D0 U1294 ( .A(n812), .B(n811), .C(n865), .ZN(n863) );
  MAOI222D0 U1295 ( .A(n863), .B(n814), .C(n813), .ZN(n859) );
  MAOI222D0 U1296 ( .A(n816), .B(n815), .C(n859), .ZN(n857) );
  MAOI222D0 U1297 ( .A(n857), .B(n818), .C(n817), .ZN(n853) );
  MAOI222D0 U1298 ( .A(n820), .B(n819), .C(n853), .ZN(n851) );
  MAOI222D0 U1299 ( .A(n851), .B(n822), .C(n821), .ZN(n847) );
  MAOI222D0 U1300 ( .A(n824), .B(n823), .C(n847), .ZN(n845) );
  MAOI222D0 U1301 ( .A(n845), .B(n826), .C(n825), .ZN(n841) );
  MAOI222D0 U1302 ( .A(n828), .B(n827), .C(n841), .ZN(n876) );
  MAOI222D0 U1303 ( .A(n876), .B(n830), .C(n829), .ZN(n872) );
  MAOI222D0 U1304 ( .A(n832), .B(n831), .C(n872), .ZN(n889) );
  MAOI222D0 U1305 ( .A(n889), .B(n834), .C(n833), .ZN(n885) );
  MAOI222D0 U1306 ( .A(n836), .B(n835), .C(n885), .ZN(n838) );
  CKND2D0 U1307 ( .A1(n838), .A2(n837), .ZN(n930) );
  OAI21D0 U1308 ( .A1(n838), .A2(n837), .B(n930), .ZN(add_tc[23]) );
  OA21D0 U1309 ( .A1(n882), .A2(n839), .B(n918), .Z(N142) );
  INVD0 U1310 ( .I(n841), .ZN(n842) );
  MUX2ND0 U1311 ( .I0(n842), .I1(n841), .S(n840), .ZN(add_tc[18]) );
  INVD0 U1312 ( .I(n845), .ZN(n844) );
  MUX2ND0 U1313 ( .I0(n845), .I1(n844), .S(n843), .ZN(add_tc[17]) );
  INVD0 U1314 ( .I(n847), .ZN(n848) );
  MUX2ND0 U1315 ( .I0(n848), .I1(n847), .S(n846), .ZN(add_tc[16]) );
  INVD0 U1316 ( .I(n851), .ZN(n850) );
  MUX2ND0 U1317 ( .I0(n851), .I1(n850), .S(n849), .ZN(add_tc[15]) );
  INVD0 U1318 ( .I(n853), .ZN(n854) );
  MUX2ND0 U1319 ( .I0(n854), .I1(n853), .S(n852), .ZN(add_tc[14]) );
  INVD0 U1320 ( .I(n857), .ZN(n856) );
  MUX2ND0 U1321 ( .I0(n857), .I1(n856), .S(n855), .ZN(add_tc[13]) );
  MUX2ND0 U1322 ( .I0(n860), .I1(n859), .S(n858), .ZN(add_tc[12]) );
  MUX2ND0 U1323 ( .I0(n863), .I1(n862), .S(n861), .ZN(add_tc[11]) );
  INVD0 U1324 ( .I(n865), .ZN(n866) );
  MUX2ND0 U1325 ( .I0(n866), .I1(n865), .S(n864), .ZN(add_tc[10]) );
  INVD0 U1326 ( .I(add_tc[17]), .ZN(n898) );
  INVD0 U1327 ( .I(add_tc[15]), .ZN(n881) );
  INVD0 U1328 ( .I(add_tc[13]), .ZN(n868) );
  INVD0 U1329 ( .I(add_tc[11]), .ZN(n926) );
  NR2D0 U1330 ( .A1(add_tc[10]), .A2(n878), .ZN(n925) );
  CKND2D0 U1331 ( .A1(n926), .A2(n925), .ZN(n924) );
  NR2D0 U1332 ( .A1(add_tc[12]), .A2(n924), .ZN(n910) );
  CKND2D0 U1333 ( .A1(n868), .A2(n910), .ZN(n877) );
  NR2D0 U1334 ( .A1(add_tc[14]), .A2(n877), .ZN(n880) );
  CKND2D0 U1335 ( .A1(n881), .A2(n880), .ZN(n879) );
  NR2D0 U1336 ( .A1(add_tc[16]), .A2(n879), .ZN(n897) );
  CKND2D0 U1337 ( .A1(n898), .A2(n897), .ZN(n896) );
  NR2D0 U1338 ( .A1(add_tc[18]), .A2(n896), .ZN(n891) );
  AOI21D0 U1339 ( .A1(add_tc[18]), .A2(n896), .B(n891), .ZN(N92) );
  AOI21D0 U1340 ( .A1(sub_tc[6]), .A2(n905), .B(n867), .ZN(N131) );
  AOI21D0 U1341 ( .A1(sub_tc[20]), .A2(n903), .B(n895), .ZN(N145) );
  OA21D0 U1342 ( .A1(n870), .A2(n869), .B(n900), .Z(N134) );
  AOI21D0 U1343 ( .A1(add_tc[6]), .A2(n901), .B(n909), .ZN(N80) );
  INVD0 U1344 ( .I(n872), .ZN(n873) );
  MUX2ND0 U1345 ( .I0(n873), .I1(n872), .S(n871), .ZN(add_tc[20]) );
  INVD0 U1346 ( .I(n876), .ZN(n875) );
  MUX2ND0 U1347 ( .I0(n876), .I1(n875), .S(n874), .ZN(add_tc[19]) );
  INVD0 U1348 ( .I(add_tc[19]), .ZN(n892) );
  CKND2D0 U1349 ( .A1(n892), .A2(n891), .ZN(n890) );
  NR2D0 U1350 ( .A1(add_tc[20]), .A2(n890), .ZN(n915) );
  AOI21D0 U1351 ( .A1(add_tc[20]), .A2(n890), .B(n915), .ZN(N94) );
  AOI21D0 U1352 ( .A1(add_tc[16]), .A2(n879), .B(n897), .ZN(N90) );
  AOI21D0 U1353 ( .A1(add_tc[14]), .A2(n877), .B(n880), .ZN(N88) );
  AOI21D0 U1354 ( .A1(add_tc[10]), .A2(n878), .B(n925), .ZN(N84) );
  OA21D0 U1355 ( .A1(n881), .A2(n880), .B(n879), .Z(N89) );
  AOI21D0 U1356 ( .A1(sub_tc[16]), .A2(n883), .B(n882), .ZN(N141) );
  INVD0 U1357 ( .I(n885), .ZN(n886) );
  MUX2ND0 U1358 ( .I0(n886), .I1(n885), .S(n884), .ZN(add_tc[22]) );
  MUX2ND0 U1359 ( .I0(n889), .I1(n888), .S(n887), .ZN(add_tc[21]) );
  INVD0 U1360 ( .I(add_tc[21]), .ZN(n916) );
  CKND2D0 U1361 ( .A1(n916), .A2(n915), .ZN(n914) );
  NR2D0 U1362 ( .A1(add_tc[22]), .A2(n914), .ZN(n2262) );
  AOI21D0 U1363 ( .A1(add_tc[22]), .A2(n914), .B(n2262), .ZN(N96) );
  OA21D0 U1364 ( .A1(n892), .A2(n891), .B(n890), .Z(N93) );
  OA21D0 U1365 ( .A1(n895), .A2(n894), .B(n893), .Z(N146) );
  OA21D0 U1366 ( .A1(n898), .A2(n897), .B(n896), .Z(N91) );
  AOI21D0 U1367 ( .A1(sub_tc[10]), .A2(n900), .B(n899), .ZN(N135) );
  OA21D0 U1368 ( .A1(n922), .A2(n902), .B(n901), .Z(N79) );
  OA21D0 U1369 ( .A1(n917), .A2(n904), .B(n903), .Z(N144) );
  OA21D0 U1370 ( .A1(n906), .A2(n912), .B(n905), .Z(N130) );
  OA21D0 U1371 ( .A1(n909), .A2(n908), .B(n907), .Z(N81) );
  AOI21D0 U1372 ( .A1(add_tc[12]), .A2(n924), .B(n910), .ZN(N86) );
  OA21D0 U1373 ( .A1(n911), .A2(n913), .B(n923), .Z(N77) );
  AOI21D0 U1374 ( .A1(add_tc[2]), .A2(n919), .B(n913), .ZN(N76) );
  OA21D0 U1375 ( .A1(n916), .A2(n915), .B(n914), .Z(N95) );
  AOI21D0 U1376 ( .A1(sub_tc[18]), .A2(n918), .B(n917), .ZN(N143) );
  OA21D0 U1377 ( .A1(n921), .A2(n920), .B(n919), .Z(N75) );
  AOI21D0 U1378 ( .A1(add_tc[4]), .A2(n923), .B(n922), .ZN(N78) );
  OA21D0 U1379 ( .A1(n926), .A2(n925), .B(n924), .Z(N85) );
  OA21D0 U1380 ( .A1(n929), .A2(n928), .B(n927), .Z(N128) );
  OAI21D0 U1381 ( .A1(n932), .A2(n931), .B(n930), .ZN(\add_sm[23] ) );
  INVD0 U1382 ( .I(\add_sm[23] ), .ZN(n70) );
  NR2D0 U1383 ( .A1(n933), .A2(n932), .ZN(n935) );
  NR2D0 U1384 ( .A1(n935), .A2(n934), .ZN(\sub_sm[23] ) );
  INVD0 U1385 ( .I(\sub_sm[23] ), .ZN(n69) );
  FA1D0 U1386 ( .A(S[16]), .B(S[17]), .CI(n936), .CO(n961), .S(n1770) );
  NR2D0 U1387 ( .A1(n1767), .A2(n1470), .ZN(n938) );
  OAI22D0 U1388 ( .A1(n1772), .A2(n1472), .B1(n1777), .B2(n1471), .ZN(n937) );
  AOI211D0 U1389 ( .A1(n1475), .A2(n1770), .B(n938), .C(n937), .ZN(n939) );
  MUX2ND0 U1390 ( .I0(n1477), .I1(R[20]), .S(n939), .ZN(n948) );
  FA1D0 U1391 ( .A(S[13]), .B(S[14]), .CI(n940), .CO(n943), .S(n1785) );
  NR2D0 U1392 ( .A1(n1782), .A2(n1417), .ZN(n942) );
  AOI211D0 U1393 ( .A1(n1385), .A2(n1785), .B(n942), .C(n941), .ZN(n947) );
  FA1D0 U1394 ( .A(S[14]), .B(S[15]), .CI(n943), .CO(n1128), .S(n1780) );
  OAI22D0 U1395 ( .A1(n1782), .A2(n1419), .B1(n1787), .B2(n1394), .ZN(n944) );
  AOI211D0 U1396 ( .A1(n1385), .A2(n1780), .B(n945), .C(n944), .ZN(n950) );
  INVD0 U1397 ( .I(n946), .ZN(\mult_x_9/n201 ) );
  FA1D0 U1398 ( .A(\mult_x_9/n203 ), .B(n948), .CI(n947), .CO(n951), .S(n949)
         );
  INVD0 U1399 ( .I(n949), .ZN(\mult_x_9/n209 ) );
  FA1D0 U1400 ( .A(\mult_x_9/n203 ), .B(n951), .CI(n950), .CO(n946), .S(n952)
         );
  INVD0 U1401 ( .I(n952), .ZN(\mult_x_9/n202 ) );
  INVD0 U1402 ( .I(inv_Q_mag[17]), .ZN(n2111) );
  NR2D0 U1403 ( .A1(n2111), .A2(n1893), .ZN(n954) );
  INVD0 U1404 ( .I(inv_Q_mag[16]), .ZN(n2115) );
  INVD0 U1405 ( .I(inv_Q_mag[15]), .ZN(n2119) );
  OAI22D0 U1406 ( .A1(n2115), .A2(n1895), .B1(n2119), .B2(n1894), .ZN(n953) );
  AOI211D0 U1407 ( .A1(n1898), .A2(n2210), .B(n954), .C(n953), .ZN(n955) );
  MUX2ND0 U1408 ( .I0(n1900), .I1(R_lat_mag[20]), .S(n955), .ZN(n965) );
  INVD0 U1409 ( .I(inv_Q_mag[12]), .ZN(n2131) );
  NR2D0 U1410 ( .A1(n2131), .A2(n1285), .ZN(n957) );
  INVD0 U1411 ( .I(inv_Q_mag[14]), .ZN(n2123) );
  OAI22D0 U1412 ( .A1(n2123), .A2(n1840), .B1(n2127), .B2(n1842), .ZN(n956) );
  AOI211D0 U1413 ( .A1(n1334), .A2(n2222), .B(n957), .C(n956), .ZN(n964) );
  OAI22D0 U1414 ( .A1(n2119), .A2(n1840), .B1(n2123), .B2(n1842), .ZN(n958) );
  AOI211D0 U1415 ( .A1(n1334), .A2(n2218), .B(n959), .C(n958), .ZN(n983) );
  INVD0 U1416 ( .I(n960), .ZN(\mult_x_13/n201 ) );
  AOI22D0 U1417 ( .A1(S[17]), .A2(n1384), .B1(S[16]), .B2(n1383), .ZN(n963) );
  FA1D0 U1418 ( .A(S[17]), .B(S[18]), .CI(n961), .CO(n1023), .S(n1765) );
  CKND2D0 U1419 ( .A1(n1765), .A2(n1385), .ZN(n962) );
  FA1D0 U1420 ( .A(\mult_x_13/n203 ), .B(n965), .CI(n964), .CO(n984), .S(n966)
         );
  INVD0 U1421 ( .I(n966), .ZN(\mult_x_13/n209 ) );
  NR2D0 U1422 ( .A1(n2131), .A2(n1893), .ZN(n968) );
  INVD0 U1423 ( .I(inv_Q_mag[10]), .ZN(n2139) );
  INVD0 U1424 ( .I(inv_Q_mag[11]), .ZN(n2135) );
  OAI22D0 U1425 ( .A1(n2139), .A2(n1894), .B1(n2135), .B2(n1895), .ZN(n967) );
  AOI211D0 U1426 ( .A1(n1898), .A2(n2230), .B(n968), .C(n967), .ZN(n969) );
  MUX2ND0 U1427 ( .I0(n1900), .I1(R_lat_mag[20]), .S(n969), .ZN(n1003) );
  NR2D0 U1428 ( .A1(n2151), .A2(n1285), .ZN(n971) );
  INVD0 U1429 ( .I(inv_Q_mag[8]), .ZN(n2147) );
  OAI22D0 U1430 ( .A1(n2147), .A2(n1842), .B1(n2143), .B2(n1840), .ZN(n970) );
  AOI211D0 U1431 ( .A1(n1334), .A2(n2242), .B(n971), .C(n970), .ZN(n1002) );
  INVD0 U1432 ( .I(n972), .ZN(\mult_x_13/n245 ) );
  FA1D0 U1433 ( .A(S[11]), .B(S[12]), .CI(n973), .CO(n575), .S(n1795) );
  NR2D0 U1434 ( .A1(n1792), .A2(n1470), .ZN(n975) );
  OAI22D0 U1435 ( .A1(n1797), .A2(n1472), .B1(n1802), .B2(n1471), .ZN(n974) );
  AOI211D0 U1436 ( .A1(n1475), .A2(n1795), .B(n975), .C(n974), .ZN(n976) );
  MUX2ND0 U1437 ( .I0(n1477), .I1(R[20]), .S(n976), .ZN(n998) );
  FA1D0 U1438 ( .A(S[8]), .B(S[9]), .CI(n977), .CO(n1099), .S(n1810) );
  NR2D0 U1439 ( .A1(n1807), .A2(n1417), .ZN(n979) );
  OAI22D0 U1440 ( .A1(n1812), .A2(n1419), .B1(n1817), .B2(n1394), .ZN(n978) );
  AOI211D0 U1441 ( .A1(n1385), .A2(n1810), .B(n979), .C(n978), .ZN(n997) );
  INVD0 U1442 ( .I(n980), .ZN(\mult_x_9/n245 ) );
  AOI22D0 U1443 ( .A1(S[3]), .A2(n1384), .B1(S[2]), .B2(n1383), .ZN(n982) );
  CKND2D0 U1444 ( .A1(n1723), .A2(n1385), .ZN(n981) );
  FA1D0 U1445 ( .A(\mult_x_13/n203 ), .B(n984), .CI(n983), .CO(n960), .S(n985)
         );
  INVD0 U1446 ( .I(n985), .ZN(\mult_x_13/n202 ) );
  AOI22D0 U1447 ( .A1(inv_Q_mag[17]), .A2(n1336), .B1(inv_Q_mag[16]), .B2(
        n1337), .ZN(n987) );
  CKND2D0 U1448 ( .A1(n2206), .A2(n1334), .ZN(n986) );
  OAI211D0 U1449 ( .A1(n1840), .A2(n2107), .B(n987), .C(n986), .ZN(
        \mult_x_13/n512 ) );
  AOI22D0 U1450 ( .A1(S[5]), .A2(n1384), .B1(S[4]), .B2(n1383), .ZN(n990) );
  FA1D0 U1451 ( .A(S[5]), .B(S[6]), .CI(n988), .CO(n578), .S(n1831) );
  OAI211D0 U1452 ( .A1(n1417), .A2(n1823), .B(n990), .C(n989), .ZN(
        \mult_x_9/n523 ) );
  INVD0 U1453 ( .I(inv_Q_mag[5]), .ZN(n2159) );
  AOI22D0 U1454 ( .A1(inv_Q_mag[4]), .A2(n1336), .B1(n2162), .B2(n1334), .ZN(
        n992) );
  CKND2D0 U1455 ( .A1(inv_Q_mag[3]), .A2(n1337), .ZN(n991) );
  OAI211D0 U1456 ( .A1(n1840), .A2(n2159), .B(n992), .C(n991), .ZN(
        \mult_x_13/n524 ) );
  AOI22D0 U1457 ( .A1(S[4]), .A2(n1384), .B1(S[3]), .B2(n1383), .ZN(n994) );
  CKND2D0 U1458 ( .A1(n1719), .A2(n1385), .ZN(n993) );
  OAI211D0 U1459 ( .A1(n1417), .A2(n1827), .B(n994), .C(n993), .ZN(
        \mult_x_9/n524 ) );
  INVD0 U1460 ( .I(inv_Q_mag[6]), .ZN(n2155) );
  AOI22D0 U1461 ( .A1(inv_Q_mag[5]), .A2(n1336), .B1(n2254), .B2(n1334), .ZN(
        n996) );
  CKND2D0 U1462 ( .A1(inv_Q_mag[4]), .A2(n1337), .ZN(n995) );
  OAI211D0 U1463 ( .A1(n1840), .A2(n2155), .B(n996), .C(n995), .ZN(
        \mult_x_13/n523 ) );
  FA1D0 U1464 ( .A(\mult_x_9/n247 ), .B(n998), .CI(n997), .CO(n980), .S(n999)
         );
  INVD0 U1465 ( .I(n999), .ZN(\mult_x_9/n246 ) );
  CKND2D0 U1466 ( .A1(n1795), .A2(n1385), .ZN(n1000) );
  OAI211D0 U1467 ( .A1(n1417), .A2(n1792), .B(n1001), .C(n1000), .ZN(
        \mult_x_9/n518 ) );
  FA1D0 U1468 ( .A(\mult_x_13/n247 ), .B(n1003), .CI(n1002), .CO(n972), .S(
        n1004) );
  INVD0 U1469 ( .I(n1004), .ZN(\mult_x_13/n246 ) );
  AOI22D0 U1470 ( .A1(inv_Q_mag[11]), .A2(n1336), .B1(n2230), .B2(n1334), .ZN(
        n1006) );
  CKND2D0 U1471 ( .A1(inv_Q_mag[10]), .A2(n1337), .ZN(n1005) );
  OAI211D0 U1472 ( .A1(n1840), .A2(n2131), .B(n1006), .C(n1005), .ZN(
        \mult_x_13/n518 ) );
  FA1D0 U1473 ( .A(S[10]), .B(S[11]), .CI(n1007), .CO(n973), .S(n1800) );
  OAI22D0 U1474 ( .A1(n1802), .A2(n1472), .B1(n1807), .B2(n1471), .ZN(n1008)
         );
  AOI211D0 U1475 ( .A1(n1475), .A2(n1800), .B(n1009), .C(n1008), .ZN(n1010) );
  MUX2ND0 U1476 ( .I0(n1477), .I1(R[20]), .S(n1010), .ZN(n1309) );
  FA1D0 U1477 ( .A(S[7]), .B(S[8]), .CI(n1011), .CO(n977), .S(n1815) );
  OAI22D0 U1478 ( .A1(n1817), .A2(n1419), .B1(n1823), .B2(n1394), .ZN(n1012)
         );
  AOI211D0 U1479 ( .A1(n1385), .A2(n1815), .B(n1013), .C(n1012), .ZN(n1308) );
  INVD0 U1480 ( .I(inv_Q_mag[4]), .ZN(n2164) );
  AOI22D0 U1481 ( .A1(inv_Q_mag[3]), .A2(n1336), .B1(n2167), .B2(n1334), .ZN(
        n1016) );
  CKND2D0 U1482 ( .A1(inv_Q_mag[2]), .A2(n1337), .ZN(n1015) );
  OAI211D0 U1483 ( .A1(n1840), .A2(n2164), .B(n1016), .C(n1015), .ZN(
        \mult_x_13/n525 ) );
  NR2D0 U1484 ( .A1(n2135), .A2(n1893), .ZN(n1018) );
  OAI22D0 U1485 ( .A1(n2143), .A2(n1894), .B1(n2139), .B2(n1895), .ZN(n1017)
         );
  AOI211D0 U1486 ( .A1(n1898), .A2(n2234), .B(n1018), .C(n1017), .ZN(n1019) );
  MUX2ND0 U1487 ( .I0(n1900), .I1(R_lat_mag[20]), .S(n1019), .ZN(n1298) );
  NR2D0 U1488 ( .A1(n2155), .A2(n1285), .ZN(n1021) );
  OAI22D0 U1489 ( .A1(n2151), .A2(n1842), .B1(n2147), .B2(n1840), .ZN(n1020)
         );
  AOI211D0 U1490 ( .A1(n1334), .A2(n2246), .B(n1021), .C(n1020), .ZN(n1297) );
  INVD0 U1491 ( .I(n1022), .ZN(\mult_x_13/n256 ) );
  FA1D0 U1492 ( .A(S[18]), .B(S[19]), .CI(n1023), .CO(n1034), .S(n1760) );
  CKND2D0 U1493 ( .A1(S[22]), .A2(n1024), .ZN(n1737) );
  OAI21D0 U1494 ( .A1(S[22]), .A2(n1024), .B(n1737), .ZN(n1739) );
  OAI222D0 U1495 ( .A1(n1394), .A2(n1747), .B1(n1419), .B2(n1742), .C1(n1421), 
        .C2(n1739), .ZN(n1396) );
  INVD0 U1496 ( .I(\mult_x_9/n178 ), .ZN(n1161) );
  FA1D0 U1497 ( .A(S[21]), .B(S[22]), .CI(n1025), .CO(n1024), .S(n1745) );
  NR2D0 U1498 ( .A1(n1742), .A2(n1417), .ZN(n1027) );
  AOI211D0 U1499 ( .A1(n1385), .A2(n1745), .B(n1027), .C(n1026), .ZN(n1160) );
  FA1D0 U1500 ( .A(S[20]), .B(S[21]), .CI(n1028), .CO(n1025), .S(n1750) );
  NR2D0 U1501 ( .A1(n1747), .A2(n1417), .ZN(n1030) );
  OAI22D0 U1502 ( .A1(n1752), .A2(n1419), .B1(n1757), .B2(n1394), .ZN(n1029)
         );
  AOI211D0 U1503 ( .A1(n1385), .A2(n1750), .B(n1030), .C(n1029), .ZN(n1033) );
  OAI22D0 U1504 ( .A1(n1742), .A2(n1471), .B1(n1037), .B2(n1737), .ZN(n1031)
         );
  MUX2ND0 U1505 ( .I0(R[20]), .I1(n1477), .S(n1031), .ZN(n1032) );
  FA1D0 U1506 ( .A(\mult_x_9/n178 ), .B(n1033), .CI(n1032), .CO(n1165), .S(
        n1169) );
  FA1D0 U1507 ( .A(S[19]), .B(S[20]), .CI(n1034), .CO(n1028), .S(n1755) );
  NR2D0 U1508 ( .A1(n1752), .A2(n1417), .ZN(n1036) );
  OAI222D0 U1509 ( .A1(n1739), .A2(n1037), .B1(n1472), .B2(n1742), .C1(n1471), 
        .C2(n1747), .ZN(n1038) );
  MUX2ND0 U1510 ( .I0(R[20]), .I1(n1477), .S(n1038), .ZN(n1158) );
  INVD0 U1511 ( .I(\mult_x_9/n186 ), .ZN(n1177) );
  INVD0 U1512 ( .I(\mult_x_9/n187 ), .ZN(n1281) );
  INVD0 U1513 ( .I(\mult_x_9/n195 ), .ZN(n1273) );
  INVD0 U1514 ( .I(\mult_x_9/n192 ), .ZN(n1272) );
  INVD0 U1515 ( .I(\mult_x_9/n199 ), .ZN(n1173) );
  INVD0 U1516 ( .I(\mult_x_9/n196 ), .ZN(n1172) );
  INVD0 U1517 ( .I(\mult_x_9/n200 ), .ZN(n1189) );
  INVD0 U1518 ( .I(\mult_x_9/n206 ), .ZN(n1188) );
  INVD0 U1519 ( .I(\mult_x_9/n212 ), .ZN(n1181) );
  INVD0 U1520 ( .I(\mult_x_9/n207 ), .ZN(n1180) );
  INVD0 U1521 ( .I(\mult_x_9/n217 ), .ZN(n1185) );
  INVD0 U1522 ( .I(\mult_x_9/n213 ), .ZN(n1184) );
  INVD0 U1523 ( .I(\mult_x_9/n218 ), .ZN(n1197) );
  INVD0 U1524 ( .I(\mult_x_9/n232 ), .ZN(n1221) );
  INVD0 U1525 ( .I(\mult_x_9/n226 ), .ZN(n1220) );
  INVD0 U1526 ( .I(\mult_x_9/n240 ), .ZN(n1265) );
  INVD0 U1527 ( .I(\mult_x_9/n233 ), .ZN(n1264) );
  INVD0 U1528 ( .I(\mult_x_9/n241 ), .ZN(n1269) );
  INVD0 U1529 ( .I(\mult_x_9/n259 ), .ZN(n1257) );
  INVD0 U1530 ( .I(\mult_x_9/n251 ), .ZN(n1256) );
  INVD0 U1531 ( .I(\mult_x_9/n267 ), .ZN(n1229) );
  INVD0 U1532 ( .I(\mult_x_9/n260 ), .ZN(n1228) );
  INVD0 U1533 ( .I(\mult_x_9/n268 ), .ZN(n1217) );
  INVD0 U1534 ( .I(\mult_x_9/n285 ), .ZN(n1237) );
  INVD0 U1535 ( .I(\mult_x_9/n277 ), .ZN(n1236) );
  INVD0 U1536 ( .I(\mult_x_9/n294 ), .ZN(n1225) );
  INVD0 U1537 ( .I(\mult_x_9/n286 ), .ZN(n1224) );
  INVD0 U1538 ( .I(\mult_x_9/n295 ), .ZN(n1205) );
  INVD0 U1539 ( .I(\mult_x_9/n304 ), .ZN(n1209) );
  INVD0 U1540 ( .I(\mult_x_9/n313 ), .ZN(n1233) );
  INVD0 U1541 ( .I(\mult_x_9/n331 ), .ZN(n1253) );
  INVD0 U1542 ( .I(\mult_x_9/n341 ), .ZN(n1241) );
  INVD0 U1543 ( .I(\mult_x_9/n361 ), .ZN(n1261) );
  INVD0 U1544 ( .I(\mult_x_9/n369 ), .ZN(n1245) );
  INVD0 U1545 ( .I(\mult_x_9/n385 ), .ZN(n1193) );
  XOR3D0 U1546 ( .A1(n1041), .A2(n1040), .A3(n1039), .Z(n1074) );
  CKXOR2D0 U1547 ( .A1(n1043), .A2(n1042), .Z(n1068) );
  AOI22D0 U1548 ( .A1(R[2]), .A2(n1044), .B1(R[1]), .B2(\mult_x_9/n686 ), .ZN(
        n1045) );
  NR2D0 U1549 ( .A1(n1046), .A2(n1045), .ZN(n1157) );
  CKND2D0 U1550 ( .A1(R[0]), .A2(n1045), .ZN(n1147) );
  NR2D0 U1551 ( .A1(n1825), .A2(n1147), .ZN(n1049) );
  CKND2D0 U1552 ( .A1(R[1]), .A2(n1046), .ZN(n1151) );
  CKND2D0 U1553 ( .A1(R[2]), .A2(n1047), .ZN(n1153) );
  OAI22D0 U1554 ( .A1(n1730), .A2(n1151), .B1(n1726), .B2(n1153), .ZN(n1048)
         );
  AOI211D0 U1555 ( .A1(n1157), .A2(n1723), .B(n1049), .C(n1048), .ZN(n1050) );
  MUX2ND0 U1556 ( .I0(\mult_x_9/n686 ), .I1(R[2]), .S(n1050), .ZN(n1062) );
  INVD0 U1557 ( .I(n1059), .ZN(n1052) );
  OAI21D0 U1558 ( .A1(n1052), .A2(\mult_x_9/n660 ), .B(n80), .ZN(n1051) );
  OAI31D0 U1559 ( .A1(n1052), .A2(n80), .A3(\mult_x_9/n660 ), .B(n1051), .ZN(
        n1061) );
  NR2D0 U1560 ( .A1(\mult_x_9/n686 ), .A2(n1053), .ZN(n1058) );
  NR2D0 U1561 ( .A1(n1730), .A2(n1147), .ZN(n1055) );
  CKND2D0 U1562 ( .A1(\mult_x_9/n686 ), .A2(n1057), .ZN(n1056) );
  OAI221D0 U1563 ( .A1(n1059), .A2(n1058), .B1(\mult_x_9/n686 ), .B2(n1057), 
        .C(n1056), .ZN(n1060) );
  MAOI222D0 U1564 ( .A(n1062), .B(n1061), .C(n1060), .ZN(n1067) );
  NR2D0 U1565 ( .A1(n1827), .A2(n1147), .ZN(n1064) );
  AOI211D0 U1566 ( .A1(n1157), .A2(n1719), .B(n1064), .C(n1063), .ZN(n1065) );
  MUX2ND0 U1567 ( .I0(R[2]), .I1(\mult_x_9/n686 ), .S(n1065), .ZN(n1066) );
  MAOI222D0 U1568 ( .A(n1068), .B(n1067), .C(n1066), .ZN(n1073) );
  NR2D0 U1569 ( .A1(n1823), .A2(n1147), .ZN(n1070) );
  OAI22D0 U1570 ( .A1(n1827), .A2(n1151), .B1(n1825), .B2(n1153), .ZN(n1069)
         );
  AOI211D0 U1571 ( .A1(n1157), .A2(n1831), .B(n1070), .C(n1069), .ZN(n1071) );
  MUX2ND0 U1572 ( .I0(\mult_x_9/n686 ), .I1(R[2]), .S(n1071), .ZN(n1072) );
  MAOI222D0 U1573 ( .A(n1074), .B(n1073), .C(n1072), .ZN(n1084) );
  NR2D0 U1574 ( .A1(n1817), .A2(n1147), .ZN(n1076) );
  OAI22D0 U1575 ( .A1(n1823), .A2(n1151), .B1(n1827), .B2(n1153), .ZN(n1075)
         );
  AOI211D0 U1576 ( .A1(n1157), .A2(n1820), .B(n1076), .C(n1075), .ZN(n1077) );
  MUX2ND0 U1577 ( .I0(R[2]), .I1(\mult_x_9/n686 ), .S(n1077), .ZN(n1083) );
  FA1D0 U1578 ( .A(n1080), .B(n1079), .CI(n1078), .CO(n1086), .S(n1081) );
  INVD0 U1579 ( .I(n1081), .ZN(n1082) );
  MAOI222D0 U1580 ( .A(n1084), .B(n1083), .C(n1082), .ZN(n1093) );
  FA1D0 U1581 ( .A(n1087), .B(n1086), .CI(n1085), .CO(n536), .S(n1092) );
  NR2D0 U1582 ( .A1(n1812), .A2(n1147), .ZN(n1089) );
  MUX2ND0 U1583 ( .I0(\mult_x_9/n686 ), .I1(R[2]), .S(n1090), .ZN(n1091) );
  MAOI222D0 U1584 ( .A(n1093), .B(n1092), .C(n1091), .ZN(n1098) );
  NR2D0 U1585 ( .A1(n1807), .A2(n1147), .ZN(n1095) );
  OAI22D0 U1586 ( .A1(n1812), .A2(n1151), .B1(n1817), .B2(n1153), .ZN(n1094)
         );
  AOI211D0 U1587 ( .A1(n1157), .A2(n1810), .B(n1095), .C(n1094), .ZN(n1096) );
  MUX2ND0 U1588 ( .I0(R[2]), .I1(\mult_x_9/n686 ), .S(n1096), .ZN(n1097) );
  MAOI222D0 U1589 ( .A(\mult_x_9/n416 ), .B(n1098), .C(n1097), .ZN(n1105) );
  FA1D0 U1590 ( .A(S[9]), .B(S[10]), .CI(n1099), .CO(n1007), .S(n1805) );
  NR2D0 U1591 ( .A1(n1802), .A2(n1147), .ZN(n1101) );
  OAI22D0 U1592 ( .A1(n1807), .A2(n1151), .B1(n1812), .B2(n1153), .ZN(n1100)
         );
  AOI211D0 U1593 ( .A1(n1157), .A2(n1805), .B(n1101), .C(n1100), .ZN(n1102) );
  MUX2ND0 U1594 ( .I0(\mult_x_9/n686 ), .I1(R[2]), .S(n1102), .ZN(n1104) );
  MAOI222D0 U1595 ( .A(n1105), .B(n1104), .C(n1103), .ZN(n1110) );
  NR2D0 U1596 ( .A1(n1797), .A2(n1147), .ZN(n1107) );
  OAI22D0 U1597 ( .A1(n1802), .A2(n1151), .B1(n1807), .B2(n1153), .ZN(n1106)
         );
  AOI211D0 U1598 ( .A1(n1157), .A2(n1800), .B(n1107), .C(n1106), .ZN(n1108) );
  MUX2ND0 U1599 ( .I0(R[2]), .I1(\mult_x_9/n686 ), .S(n1108), .ZN(n1109) );
  MAOI222D0 U1600 ( .A(\mult_x_9/n406 ), .B(n1110), .C(n1109), .ZN(n1116) );
  NR2D0 U1601 ( .A1(n1792), .A2(n1147), .ZN(n1112) );
  OAI22D0 U1602 ( .A1(n1797), .A2(n1151), .B1(n1802), .B2(n1153), .ZN(n1111)
         );
  AOI211D0 U1603 ( .A1(n1157), .A2(n1795), .B(n1112), .C(n1111), .ZN(n1113) );
  MUX2ND0 U1604 ( .I0(\mult_x_9/n686 ), .I1(R[2]), .S(n1113), .ZN(n1115) );
  INVD0 U1605 ( .I(\mult_x_9/n399 ), .ZN(n1114) );
  MAOI222D0 U1606 ( .A(n1116), .B(n1115), .C(n1114), .ZN(n1121) );
  NR2D0 U1607 ( .A1(n1787), .A2(n1147), .ZN(n1118) );
  OAI22D0 U1608 ( .A1(n1792), .A2(n1151), .B1(n1797), .B2(n1153), .ZN(n1117)
         );
  AOI211D0 U1609 ( .A1(n1157), .A2(n1790), .B(n1118), .C(n1117), .ZN(n1119) );
  MUX2ND0 U1610 ( .I0(R[2]), .I1(\mult_x_9/n686 ), .S(n1119), .ZN(n1120) );
  MAOI222D0 U1611 ( .A(\mult_x_9/n392 ), .B(n1121), .C(n1120), .ZN(n1192) );
  NR2D0 U1612 ( .A1(n1782), .A2(n1147), .ZN(n1123) );
  OAI22D0 U1613 ( .A1(n1787), .A2(n1151), .B1(n1792), .B2(n1153), .ZN(n1122)
         );
  AOI211D0 U1614 ( .A1(n1785), .A2(n1157), .B(n1123), .C(n1122), .ZN(n1124) );
  MUX2ND0 U1615 ( .I0(\mult_x_9/n686 ), .I1(R[2]), .S(n1124), .ZN(n1191) );
  NR2D0 U1616 ( .A1(n1777), .A2(n1147), .ZN(n1126) );
  OAI22D0 U1617 ( .A1(n1782), .A2(n1151), .B1(n1787), .B2(n1153), .ZN(n1125)
         );
  AOI211D0 U1618 ( .A1(n1780), .A2(n1157), .B(n1126), .C(n1125), .ZN(n1127) );
  MUX2ND0 U1619 ( .I0(\mult_x_9/n686 ), .I1(R[2]), .S(n1127), .ZN(n1211) );
  FA1D0 U1620 ( .A(S[15]), .B(S[16]), .CI(n1128), .CO(n936), .S(n1775) );
  NR2D0 U1621 ( .A1(n1772), .A2(n1147), .ZN(n1130) );
  AOI211D0 U1622 ( .A1(n1775), .A2(n1157), .B(n1130), .C(n1129), .ZN(n1131) );
  MUX2ND0 U1623 ( .I0(\mult_x_9/n686 ), .I1(R[2]), .S(n1131), .ZN(n1243) );
  NR2D0 U1624 ( .A1(n1767), .A2(n1147), .ZN(n1133) );
  OAI22D0 U1625 ( .A1(n1772), .A2(n1151), .B1(n1777), .B2(n1153), .ZN(n1132)
         );
  MUX2ND0 U1626 ( .I0(\mult_x_9/n686 ), .I1(R[2]), .S(n1134), .ZN(n1259) );
  NR2D0 U1627 ( .A1(n1762), .A2(n1147), .ZN(n1136) );
  OAI22D0 U1628 ( .A1(n1767), .A2(n1151), .B1(n1772), .B2(n1153), .ZN(n1135)
         );
  AOI211D0 U1629 ( .A1(n1765), .A2(n1157), .B(n1136), .C(n1135), .ZN(n1137) );
  MUX2ND0 U1630 ( .I0(\mult_x_9/n686 ), .I1(R[2]), .S(n1137), .ZN(n1199) );
  NR2D0 U1631 ( .A1(n1757), .A2(n1147), .ZN(n1139) );
  OAI22D0 U1632 ( .A1(n1762), .A2(n1151), .B1(n1767), .B2(n1153), .ZN(n1138)
         );
  AOI211D0 U1633 ( .A1(n1760), .A2(n1157), .B(n1139), .C(n1138), .ZN(n1140) );
  MUX2ND0 U1634 ( .I0(\mult_x_9/n686 ), .I1(R[2]), .S(n1140), .ZN(n1239) );
  NR2D0 U1635 ( .A1(n1752), .A2(n1147), .ZN(n1142) );
  OAI22D0 U1636 ( .A1(n1757), .A2(n1151), .B1(n1762), .B2(n1153), .ZN(n1141)
         );
  AOI211D0 U1637 ( .A1(n1755), .A2(n1157), .B(n1142), .C(n1141), .ZN(n1143) );
  MUX2ND0 U1638 ( .I0(\mult_x_9/n686 ), .I1(R[2]), .S(n1143), .ZN(n1251) );
  NR2D0 U1639 ( .A1(n1747), .A2(n1147), .ZN(n1145) );
  OAI22D0 U1640 ( .A1(n1752), .A2(n1151), .B1(n1757), .B2(n1153), .ZN(n1144)
         );
  AOI211D0 U1641 ( .A1(n1750), .A2(n1157), .B(n1145), .C(n1144), .ZN(n1146) );
  MUX2ND0 U1642 ( .I0(\mult_x_9/n686 ), .I1(R[2]), .S(n1146), .ZN(n1247) );
  NR2D0 U1643 ( .A1(n1742), .A2(n1147), .ZN(n1149) );
  OAI22D0 U1644 ( .A1(n1747), .A2(n1151), .B1(n1752), .B2(n1153), .ZN(n1148)
         );
  AOI211D0 U1645 ( .A1(n1745), .A2(n1157), .B(n1149), .C(n1148), .ZN(n1150) );
  MUX2ND0 U1646 ( .I0(\mult_x_9/n686 ), .I1(R[2]), .S(n1150), .ZN(n1231) );
  INVD0 U1647 ( .I(n1157), .ZN(n1154) );
  OAI222D0 U1648 ( .A1(n1153), .A2(n1747), .B1(n1151), .B2(n1742), .C1(n1154), 
        .C2(n1739), .ZN(n1152) );
  MUX2ND0 U1649 ( .I0(R[2]), .I1(\mult_x_9/n686 ), .S(n1152), .ZN(n1207) );
  INVD0 U1650 ( .I(n1737), .ZN(n1156) );
  OA22D0 U1651 ( .A1(n1154), .A2(n1737), .B1(n1742), .B2(n1153), .Z(n1155) );
  FA1D0 U1652 ( .A(\mult_x_9/n178 ), .B(n1159), .CI(n1158), .CO(n1168), .S(
        n1275) );
  FA1D0 U1653 ( .A(R[20]), .B(n1161), .CI(n1160), .CO(n1393), .S(n1163) );
  FA1D0 U1654 ( .A(n1165), .B(n1164), .CI(n1163), .CO(n1392), .S(n1166) );
  INVD0 U1655 ( .I(n1166), .ZN(prod_full[43]) );
  FA1D0 U1656 ( .A(n1169), .B(n1168), .CI(n1167), .CO(n1164), .S(n1170) );
  INVD0 U1657 ( .I(n1170), .ZN(prod_full[42]) );
  FA1D0 U1658 ( .A(n1173), .B(n1172), .CI(n1171), .CO(n1271), .S(n1174) );
  INVD0 U1659 ( .I(n1174), .ZN(prod_full[37]) );
  FA1D0 U1660 ( .A(n1177), .B(n1176), .CI(n1175), .CO(n1276), .S(n1178) );
  INVD0 U1661 ( .I(n1178), .ZN(prod_full[40]) );
  FA1D0 U1662 ( .A(n1181), .B(n1180), .CI(n1179), .CO(n1187), .S(n1182) );
  FA1D0 U1663 ( .A(n1185), .B(n1184), .CI(n1183), .CO(n1179), .S(n1186) );
  INVD0 U1664 ( .I(n1186), .ZN(prod_full[34]) );
  FA1D0 U1665 ( .A(n1189), .B(n1188), .CI(n1187), .CO(n1171), .S(n1190) );
  INVD0 U1666 ( .I(n1190), .ZN(prod_full[36]) );
  FA1D0 U1667 ( .A(n1193), .B(n1192), .CI(n1191), .CO(n1212), .S(n1194) );
  FA1D0 U1668 ( .A(n1197), .B(n1196), .CI(n1195), .CO(n1183), .S(n1198) );
  INVD0 U1669 ( .I(n1198), .ZN(prod_full[33]) );
  FA1D0 U1670 ( .A(n1201), .B(n1200), .CI(n1199), .CO(n1240), .S(n1202) );
  INVD0 U1671 ( .I(n1202), .ZN(prod_full[18]) );
  FA1D0 U1672 ( .A(n1205), .B(n1204), .CI(n1203), .CO(n1223), .S(n1206) );
  INVD0 U1673 ( .I(n1206), .ZN(prod_full[24]) );
  FA1D0 U1674 ( .A(n1209), .B(n1208), .CI(n1207), .CO(n1204), .S(n1210) );
  FA1D0 U1675 ( .A(n1213), .B(n1212), .CI(n1211), .CO(n1244), .S(n1214) );
  INVD0 U1676 ( .I(n1214), .ZN(prod_full[15]) );
  FA1D0 U1677 ( .A(n1217), .B(n1216), .CI(n1215), .CO(n1227), .S(n1218) );
  INVD0 U1678 ( .I(n1218), .ZN(prod_full[27]) );
  FA1D0 U1679 ( .A(n1221), .B(n1220), .CI(n1219), .CO(n1195), .S(n1222) );
  FA1D0 U1680 ( .A(n1225), .B(n1224), .CI(n1223), .CO(n1235), .S(n1226) );
  INVD0 U1681 ( .I(n1226), .ZN(prod_full[25]) );
  FA1D0 U1682 ( .A(n1229), .B(n1228), .CI(n1227), .CO(n1255), .S(n1230) );
  INVD0 U1683 ( .I(n1230), .ZN(prod_full[28]) );
  FA1D0 U1684 ( .A(n1233), .B(n1232), .CI(n1231), .CO(n1208), .S(n1234) );
  INVD0 U1685 ( .I(n1234), .ZN(prod_full[22]) );
  FA1D0 U1686 ( .A(n1237), .B(n1236), .CI(n1235), .CO(n1215), .S(n1238) );
  INVD0 U1687 ( .I(n1238), .ZN(prod_full[26]) );
  FA1D0 U1688 ( .A(n1241), .B(n1240), .CI(n1239), .CO(n1252), .S(n1242) );
  INVD0 U1689 ( .I(n1242), .ZN(prod_full[19]) );
  FA1D0 U1690 ( .A(n1245), .B(n1244), .CI(n1243), .CO(n1260), .S(n1246) );
  INVD0 U1691 ( .I(n1246), .ZN(prod_full[16]) );
  FA1D0 U1692 ( .A(n1249), .B(n1248), .CI(n1247), .CO(n1232), .S(n1250) );
  INVD0 U1693 ( .I(n1250), .ZN(prod_full[21]) );
  FA1D0 U1694 ( .A(n1253), .B(n1252), .CI(n1251), .CO(n1248), .S(n1254) );
  INVD0 U1695 ( .I(n1254), .ZN(prod_full[20]) );
  FA1D0 U1696 ( .A(n1257), .B(n1256), .CI(n1255), .CO(n1267), .S(n1258) );
  FA1D0 U1697 ( .A(n1261), .B(n1260), .CI(n1259), .CO(n1200), .S(n1262) );
  INVD0 U1698 ( .I(n1262), .ZN(prod_full[17]) );
  FA1D0 U1699 ( .A(n1265), .B(n1264), .CI(n1263), .CO(n1219), .S(n1266) );
  INVD0 U1700 ( .I(n1266), .ZN(prod_full[31]) );
  FA1D0 U1701 ( .A(n1269), .B(n1268), .CI(n1267), .CO(n1263), .S(n1270) );
  INVD0 U1702 ( .I(n1270), .ZN(prod_full[30]) );
  FA1D0 U1703 ( .A(n1273), .B(n1272), .CI(n1271), .CO(n1279), .S(n1274) );
  INVD0 U1704 ( .I(n1274), .ZN(prod_full[38]) );
  FA1D0 U1705 ( .A(n1277), .B(n1276), .CI(n1275), .CO(n1167), .S(n1278) );
  INVD0 U1706 ( .I(n1278), .ZN(prod_full[41]) );
  FA1D0 U1707 ( .A(n1281), .B(n1280), .CI(n1279), .CO(n1175), .S(n1282) );
  INVD0 U1708 ( .I(n1282), .ZN(prod_full[39]) );
  AOI22D0 U1709 ( .A1(inv_Q_mag[16]), .A2(n1336), .B1(inv_Q_mag[15]), .B2(
        n1337), .ZN(n1284) );
  CKND2D0 U1710 ( .A1(n2210), .A2(n1334), .ZN(n1283) );
  OAI211D0 U1711 ( .A1(n1840), .A2(n2111), .B(n1284), .C(n1283), .ZN(
        \mult_x_13/n513 ) );
  INVD0 U1712 ( .I(\mult_x_13/n247 ), .ZN(n1301) );
  NR2D0 U1713 ( .A1(n2147), .A2(n1285), .ZN(n1287) );
  OAI22D0 U1714 ( .A1(n2143), .A2(n1842), .B1(n2139), .B2(n1840), .ZN(n1286)
         );
  AOI211D0 U1715 ( .A1(n1334), .A2(n2238), .B(n1287), .C(n1286), .ZN(n1300) );
  INVD0 U1716 ( .I(n1288), .ZN(\mult_x_13/n238 ) );
  INVD0 U1717 ( .I(inv_Q_mag[3]), .ZN(n2172) );
  CKND2D0 U1718 ( .A1(inv_Q_mag[1]), .A2(n1337), .ZN(n1289) );
  AOI22D0 U1719 ( .A1(inv_Q_mag[15]), .A2(n1336), .B1(n2214), .B2(n1334), .ZN(
        n1292) );
  CKND2D0 U1720 ( .A1(inv_Q_mag[14]), .A2(n1337), .ZN(n1291) );
  OAI211D0 U1721 ( .A1(n1840), .A2(n2115), .B(n1292), .C(n1291), .ZN(n1833) );
  INVD0 U1722 ( .I(\mult_x_13/n188 ), .ZN(\mult_x_13/n193 ) );
  AOI22D0 U1723 ( .A1(S[10]), .A2(n1384), .B1(S[9]), .B2(n1383), .ZN(n1294) );
  CKND2D0 U1724 ( .A1(n1800), .A2(n1385), .ZN(n1293) );
  OAI211D0 U1725 ( .A1(n1417), .A2(n1797), .B(n1294), .C(n1293), .ZN(
        \mult_x_9/n222 ) );
  INVD0 U1726 ( .I(\mult_x_9/n222 ), .ZN(\mult_x_9/n230 ) );
  AOI22D0 U1727 ( .A1(inv_Q_mag[10]), .A2(n1336), .B1(n2234), .B2(n1334), .ZN(
        n1296) );
  CKND2D0 U1728 ( .A1(inv_Q_mag[9]), .A2(n1337), .ZN(n1295) );
  OAI211D0 U1729 ( .A1(n1840), .A2(n2135), .B(n1296), .C(n1295), .ZN(
        \mult_x_13/n222 ) );
  INVD0 U1730 ( .I(\mult_x_13/n222 ), .ZN(\mult_x_13/n230 ) );
  FA1D0 U1731 ( .A(\mult_x_13/n247 ), .B(n1298), .CI(n1297), .CO(n1299), .S(
        n1022) );
  INVD0 U1732 ( .I(n1299), .ZN(\mult_x_13/n255 ) );
  FA1D0 U1733 ( .A(R_lat_mag[8]), .B(n1301), .CI(n1300), .CO(n1302), .S(n1288)
         );
  INVD0 U1734 ( .I(n1302), .ZN(\mult_x_13/n237 ) );
  INVD0 U1735 ( .I(\mult_x_9/n247 ), .ZN(n1312) );
  NR2D0 U1736 ( .A1(n1802), .A2(n1417), .ZN(n1304) );
  OAI22D0 U1737 ( .A1(n1807), .A2(n1419), .B1(n1812), .B2(n1394), .ZN(n1303)
         );
  AOI211D0 U1738 ( .A1(n1385), .A2(n1805), .B(n1304), .C(n1303), .ZN(n1311) );
  INVD0 U1739 ( .I(n1305), .ZN(\mult_x_9/n238 ) );
  AOI22D0 U1740 ( .A1(S[2]), .A2(n1384), .B1(S[1]), .B2(n1383), .ZN(n1307) );
  CKND2D0 U1741 ( .A1(n1733), .A2(n1385), .ZN(n1306) );
  OAI211D0 U1742 ( .A1(n1417), .A2(n1730), .B(n1307), .C(n1306), .ZN(
        \mult_x_9/n526 ) );
  FA1D0 U1743 ( .A(\mult_x_9/n247 ), .B(n1309), .CI(n1308), .CO(n1310), .S(
        n1014) );
  INVD0 U1744 ( .I(n1310), .ZN(\mult_x_9/n255 ) );
  FA1D0 U1745 ( .A(R[8]), .B(n1312), .CI(n1311), .CO(n1313), .S(n1305) );
  AOI211D0 U1746 ( .A1(\mult_x_9/n556 ), .A2(n1316), .B(n1315), .C(n1314), 
        .ZN(n1317) );
  AOI211D0 U1747 ( .A1(\mult_x_13/n556 ), .A2(n1320), .B(n1319), .C(n1318), 
        .ZN(n1321) );
  NR2D0 U1748 ( .A1(n1402), .A2(n1321), .ZN(\mult_x_13/n366 ) );
  AOI22D0 U1749 ( .A1(S[0]), .A2(n1383), .B1(S[1]), .B2(n1384), .ZN(n1324) );
  CKND2D0 U1750 ( .A1(S[2]), .A2(n1322), .ZN(n1323) );
  OAI211D0 U1751 ( .A1(n1421), .A2(n1325), .B(n1324), .C(n1323), .ZN(
        \mult_x_9/n527 ) );
  FA1D0 U1752 ( .A(n1328), .B(n1327), .CI(n1326), .CO(n1341), .S(n1329) );
  INVD0 U1753 ( .I(n1329), .ZN(\mult_x_9/n346 ) );
  FA1D0 U1754 ( .A(n1332), .B(n1331), .CI(n1330), .CO(n1345), .S(n1333) );
  INVD0 U1755 ( .I(n1333), .ZN(\mult_x_13/n346 ) );
  AOI22D0 U1756 ( .A1(inv_Q_mag[1]), .A2(n1336), .B1(n1335), .B2(n1334), .ZN(
        n1339) );
  CKND2D0 U1757 ( .A1(inv_Q_mag[0]), .A2(n1337), .ZN(n1338) );
  OAI211D0 U1758 ( .A1(n1840), .A2(n2170), .B(n1339), .C(n1338), .ZN(
        \mult_x_13/n527 ) );
  FA1D0 U1759 ( .A(n1342), .B(n1341), .CI(n1340), .CO(n448), .S(n1343) );
  FA1D0 U1760 ( .A(n1346), .B(n1345), .CI(n1344), .CO(n506), .S(n1347) );
  FA1D0 U1761 ( .A(n1350), .B(n1349), .CI(n1348), .CO(n477), .S(n1351) );
  INVD0 U1762 ( .I(n1351), .ZN(\mult_x_9/n387 ) );
  AOI211D0 U1763 ( .A1(\mult_x_9/n608 ), .A2(n1354), .B(n1353), .C(n1352), 
        .ZN(n1355) );
  NR2D0 U1764 ( .A1(n1405), .A2(n1355), .ZN(\mult_x_9/n408 ) );
  FA1D0 U1765 ( .A(n1358), .B(n1357), .CI(n1356), .CO(n1349), .S(n1359) );
  FA1D0 U1766 ( .A(n1362), .B(n1361), .CI(n1360), .CO(n1369), .S(n1363) );
  AOI211D0 U1767 ( .A1(\mult_x_13/n608 ), .A2(n1366), .B(n1365), .C(n1364), 
        .ZN(n1367) );
  FA1D0 U1768 ( .A(n1370), .B(n1369), .CI(n1368), .CO(n567), .S(n1371) );
  INVD0 U1769 ( .I(n1371), .ZN(\mult_x_13/n387 ) );
  NR4D0 U1770 ( .A1(S_lat_mag[2]), .A2(S_lat_mag[22]), .A3(S_lat_mag[12]), 
        .A4(S_lat_mag[14]), .ZN(n1378) );
  NR4D0 U1771 ( .A1(S_lat_mag[10]), .A2(S_lat_mag[9]), .A3(S_lat_mag[11]), 
        .A4(S_lat_mag[7]), .ZN(n1377) );
  OR4D0 U1772 ( .A1(S_lat_mag[16]), .A2(S_lat_mag[15]), .A3(S_lat_mag[17]), 
        .A4(S_lat_mag[13]), .Z(n1375) );
  NR4D0 U1773 ( .A1(S_lat_mag[4]), .A2(S_lat_mag[3]), .A3(S_lat_mag[5]), .A4(
        S_lat_mag[1]), .ZN(n1373) );
  NR4D0 U1774 ( .A1(S_lat_mag[21]), .A2(S_lat_mag[19]), .A3(S_lat_mag[18]), 
        .A4(S_lat_mag[20]), .ZN(n1372) );
  NR4D0 U1775 ( .A1(S_lat_mag[6]), .A2(S_lat_mag[8]), .A3(n1375), .A4(n1374), 
        .ZN(n1376) );
  AO31D0 U1776 ( .A1(n1378), .A2(n1377), .A3(n1376), .B(S_lat_mag[0]), .Z(
        \S_mag_safe[0] ) );
  AOI22D0 U1777 ( .A1(S[15]), .A2(n1384), .B1(S[14]), .B2(n1383), .ZN(n1382)
         );
  CKND2D0 U1778 ( .A1(n1775), .A2(n1385), .ZN(n1381) );
  INVD0 U1779 ( .I(\mult_x_9/n188 ), .ZN(\mult_x_9/n193 ) );
  AOI22D0 U1780 ( .A1(S[16]), .A2(n1384), .B1(S[15]), .B2(n1383), .ZN(n1387)
         );
  CKND2D0 U1781 ( .A1(n1770), .A2(n1385), .ZN(n1386) );
  OAI211D0 U1782 ( .A1(n1417), .A2(n1767), .B(n1387), .C(n1386), .ZN(
        \mult_x_9/n513 ) );
  INR2D0 U1783 ( .A1(ctl_d[0]), .B1(ctl_d[1]), .ZN(n78) );
  NR2D0 U1784 ( .A1(ctl_d[1]), .A2(ctl_d[0]), .ZN(n77) );
  INR2D0 U1785 ( .A1(ctl_d[1]), .B1(ctl_d[0]), .ZN(n79) );
  AOI22D0 U1786 ( .A1(\sub_sm[23] ), .A2(n78), .B1(n77), .B2(\add_sm[23] ), 
        .ZN(n1391) );
  OAI221D0 U1787 ( .A1(R[23]), .A2(S[23]), .B1(n1389), .B2(n1388), .C(n79), 
        .ZN(n1390) );
  CKND2D0 U1788 ( .A1(n1391), .A2(n1390), .ZN(result_comb[23]) );
  ND4D0 U1789 ( .A1(n74), .A2(n63), .A3(n65), .A4(n64), .ZN(result_comb[3]) );
  ND4D0 U1790 ( .A1(n74), .A2(n60), .A3(n62), .A4(n61), .ZN(result_comb[4]) );
  ND4D0 U1791 ( .A1(n74), .A2(n66), .A3(n68), .A4(n67), .ZN(result_comb[2]) );
  ND4D0 U1792 ( .A1(n74), .A2(n54), .A3(n56), .A4(n55), .ZN(result_comb[6]) );
  ND4D0 U1793 ( .A1(n74), .A2(n51), .A3(n53), .A4(n52), .ZN(result_comb[7]) );
  CKXOR2D0 U1794 ( .A1(\S_lat[23] ), .A2(\R_lat[23] ), .Z(\div_sm[23] ) );
  FA1D0 U1795 ( .A(n1396), .B(n1393), .CI(n1392), .CO(n1397), .S(n1162) );
  OAI22D0 U1796 ( .A1(n1742), .A2(n1394), .B1(n1737), .B2(n1421), .ZN(n1395)
         );
  XOR3D0 U1797 ( .A1(n1397), .A2(n1396), .A3(n1395), .Z(prod_full[45]) );
  XOR3D0 U1798 ( .A1(n1400), .A2(n1399), .A3(n1398), .Z(\mult_x_9/n356 ) );
  XOR3D0 U1799 ( .A1(n1403), .A2(n1402), .A3(n1401), .Z(\mult_x_13/n356 ) );
  XOR3D0 U1800 ( .A1(n1406), .A2(n1405), .A3(n1404), .Z(\mult_x_9/n401 ) );
  XOR3D0 U1801 ( .A1(n1409), .A2(n1408), .A3(n1407), .Z(\mult_x_13/n401 ) );
  FA1D0 U1802 ( .A(n1603), .B(\mult_x_9/n203 ), .CI(n1410), .CO(
        \mult_x_9/n188 ), .S(\mult_x_9/n197 ) );
  INVD0 U1803 ( .I(n1413), .ZN(n1412) );
  CKND2D0 U1804 ( .A1(R[17]), .A2(\mult_x_9/n382 ), .ZN(n1411) );
  MUX2ND0 U1805 ( .I0(n1413), .I1(n1412), .S(n1411), .ZN(\mult_x_9/n374 ) );
  INVD0 U1806 ( .I(n1416), .ZN(n1415) );
  CKND2D0 U1807 ( .A1(R[11]), .A2(\mult_x_9/n418 ), .ZN(n1414) );
  MUX2ND0 U1808 ( .I0(n1416), .I1(n1415), .S(n1414), .ZN(\mult_x_9/n413 ) );
  OAI222D0 U1809 ( .A1(n1421), .A2(n1420), .B1(n1419), .B2(n1418), .C1(n1728), 
        .C2(n1417), .ZN(\mult_x_9/n528 ) );
  NR2D0 U1810 ( .A1(n1742), .A2(n1470), .ZN(n1423) );
  OAI22D0 U1811 ( .A1(n1747), .A2(n1472), .B1(n1752), .B2(n1471), .ZN(n1422)
         );
  AOI211D0 U1812 ( .A1(n1475), .A2(n1745), .B(n1423), .C(n1422), .ZN(n1424) );
  MUX2ND0 U1813 ( .I0(R[20]), .I1(n1477), .S(n1424), .ZN(\mult_x_9/n533 ) );
  NR2D0 U1814 ( .A1(n1747), .A2(n1470), .ZN(n1426) );
  OAI22D0 U1815 ( .A1(n1752), .A2(n1472), .B1(n1757), .B2(n1471), .ZN(n1425)
         );
  AOI211D0 U1816 ( .A1(n1475), .A2(n1750), .B(n1426), .C(n1425), .ZN(n1427) );
  MUX2ND0 U1817 ( .I0(R[20]), .I1(n1477), .S(n1427), .ZN(\mult_x_9/n534 ) );
  NR2D0 U1818 ( .A1(n1752), .A2(n1470), .ZN(n1429) );
  OAI22D0 U1819 ( .A1(n1757), .A2(n1472), .B1(n1762), .B2(n1471), .ZN(n1428)
         );
  AOI211D0 U1820 ( .A1(n1475), .A2(n1755), .B(n1429), .C(n1428), .ZN(n1430) );
  MUX2ND0 U1821 ( .I0(R[20]), .I1(n1477), .S(n1430), .ZN(\mult_x_9/n535 ) );
  NR2D0 U1822 ( .A1(n1757), .A2(n1470), .ZN(n1432) );
  AOI211D0 U1823 ( .A1(n1475), .A2(n1760), .B(n1432), .C(n1431), .ZN(n1433) );
  MUX2ND0 U1824 ( .I0(R[20]), .I1(n1477), .S(n1433), .ZN(\mult_x_9/n536 ) );
  NR2D0 U1825 ( .A1(n1762), .A2(n1470), .ZN(n1435) );
  OAI22D0 U1826 ( .A1(n1767), .A2(n1472), .B1(n1772), .B2(n1471), .ZN(n1434)
         );
  AOI211D0 U1827 ( .A1(n1475), .A2(n1765), .B(n1435), .C(n1434), .ZN(n1436) );
  MUX2ND0 U1828 ( .I0(R[20]), .I1(n1477), .S(n1436), .ZN(\mult_x_9/n537 ) );
  NR2D0 U1829 ( .A1(n1772), .A2(n1470), .ZN(n1438) );
  OAI22D0 U1830 ( .A1(n1777), .A2(n1472), .B1(n1782), .B2(n1471), .ZN(n1437)
         );
  AOI211D0 U1831 ( .A1(n1475), .A2(n1775), .B(n1438), .C(n1437), .ZN(n1439) );
  MUX2ND0 U1832 ( .I0(R[20]), .I1(n1477), .S(n1439), .ZN(\mult_x_9/n539 ) );
  NR2D0 U1833 ( .A1(n1782), .A2(n1472), .ZN(n1441) );
  OAI22D0 U1834 ( .A1(n1777), .A2(n1470), .B1(n1787), .B2(n1471), .ZN(n1440)
         );
  AOI211D0 U1835 ( .A1(n1475), .A2(n1780), .B(n1441), .C(n1440), .ZN(n1442) );
  MUX2ND0 U1836 ( .I0(R[20]), .I1(n1477), .S(n1442), .ZN(\mult_x_9/n540 ) );
  OAI22D0 U1837 ( .A1(n1782), .A2(n1470), .B1(n1792), .B2(n1471), .ZN(n1443)
         );
  AOI211D0 U1838 ( .A1(n1475), .A2(n1785), .B(n1444), .C(n1443), .ZN(n1445) );
  MUX2ND0 U1839 ( .I0(R[20]), .I1(n1477), .S(n1445), .ZN(\mult_x_9/n541 ) );
  NR2D0 U1840 ( .A1(n1787), .A2(n1470), .ZN(n1447) );
  OAI22D0 U1841 ( .A1(n1792), .A2(n1472), .B1(n1797), .B2(n1471), .ZN(n1446)
         );
  AOI211D0 U1842 ( .A1(n1475), .A2(n1790), .B(n1447), .C(n1446), .ZN(n1448) );
  MUX2ND0 U1843 ( .I0(R[20]), .I1(n1477), .S(n1448), .ZN(\mult_x_9/n542 ) );
  NR2D0 U1844 ( .A1(n1802), .A2(n1470), .ZN(n1450) );
  OAI22D0 U1845 ( .A1(n1807), .A2(n1472), .B1(n1812), .B2(n1471), .ZN(n1449)
         );
  AOI211D0 U1846 ( .A1(n1475), .A2(n1805), .B(n1450), .C(n1449), .ZN(n1451) );
  MUX2ND0 U1847 ( .I0(R[20]), .I1(n1477), .S(n1451), .ZN(\mult_x_9/n545 ) );
  NR2D0 U1848 ( .A1(n1807), .A2(n1470), .ZN(n1453) );
  OAI22D0 U1849 ( .A1(n1812), .A2(n1472), .B1(n1817), .B2(n1471), .ZN(n1452)
         );
  AOI211D0 U1850 ( .A1(n1475), .A2(n1810), .B(n1453), .C(n1452), .ZN(n1454) );
  MUX2ND0 U1851 ( .I0(R[20]), .I1(n1477), .S(n1454), .ZN(\mult_x_9/n546 ) );
  NR2D0 U1852 ( .A1(n1812), .A2(n1470), .ZN(n1456) );
  OAI22D0 U1853 ( .A1(n1817), .A2(n1472), .B1(n1823), .B2(n1471), .ZN(n1455)
         );
  AOI211D0 U1854 ( .A1(n1475), .A2(n1815), .B(n1456), .C(n1455), .ZN(n1457) );
  MUX2ND0 U1855 ( .I0(R[20]), .I1(n1477), .S(n1457), .ZN(\mult_x_9/n547 ) );
  NR2D0 U1856 ( .A1(n1817), .A2(n1470), .ZN(n1459) );
  OAI22D0 U1857 ( .A1(n1823), .A2(n1472), .B1(n1827), .B2(n1471), .ZN(n1458)
         );
  AOI211D0 U1858 ( .A1(n1475), .A2(n1820), .B(n1459), .C(n1458), .ZN(n1460) );
  MUX2ND0 U1859 ( .I0(R[20]), .I1(n1477), .S(n1460), .ZN(\mult_x_9/n548 ) );
  NR2D0 U1860 ( .A1(n1823), .A2(n1470), .ZN(n1462) );
  OAI22D0 U1861 ( .A1(n1827), .A2(n1472), .B1(n1825), .B2(n1471), .ZN(n1461)
         );
  AOI211D0 U1862 ( .A1(n1475), .A2(n1831), .B(n1462), .C(n1461), .ZN(n1463) );
  MUX2ND0 U1863 ( .I0(R[20]), .I1(n1477), .S(n1463), .ZN(\mult_x_9/n549 ) );
  NR2D0 U1864 ( .A1(n1827), .A2(n1470), .ZN(n1465) );
  OAI22D0 U1865 ( .A1(n1825), .A2(n1472), .B1(n1730), .B2(n1471), .ZN(n1464)
         );
  MUX2ND0 U1866 ( .I0(R[20]), .I1(n1477), .S(n1466), .ZN(\mult_x_9/n550 ) );
  NR2D0 U1867 ( .A1(n1825), .A2(n1470), .ZN(n1468) );
  OAI22D0 U1868 ( .A1(n1730), .A2(n1472), .B1(n1726), .B2(n1471), .ZN(n1467)
         );
  AOI211D0 U1869 ( .A1(n1475), .A2(n1723), .B(n1468), .C(n1467), .ZN(n1469) );
  MUX2ND0 U1870 ( .I0(R[20]), .I1(n1477), .S(n1469), .ZN(\mult_x_9/n551 ) );
  NR2D0 U1871 ( .A1(n1730), .A2(n1470), .ZN(n1474) );
  OAI22D0 U1872 ( .A1(n1726), .A2(n1472), .B1(n1728), .B2(n1471), .ZN(n1473)
         );
  AOI211D0 U1873 ( .A1(n1475), .A2(n1733), .B(n1474), .C(n1473), .ZN(n1476) );
  MUX2ND0 U1874 ( .I0(R[20]), .I1(n1477), .S(n1476), .ZN(\mult_x_9/n552 ) );
  OAI22D0 U1875 ( .A1(n1742), .A2(n1530), .B1(n1479), .B2(n1737), .ZN(n1478)
         );
  MUX2ND0 U1876 ( .I0(\mult_x_9/n556 ), .I1(R[17]), .S(n1478), .ZN(
        \mult_x_9/n557 ) );
  OAI222D0 U1877 ( .A1(n1530), .A2(n1747), .B1(n1531), .B2(n1742), .C1(n1479), 
        .C2(n1739), .ZN(n1480) );
  MUX2ND0 U1878 ( .I0(\mult_x_9/n556 ), .I1(R[17]), .S(n1480), .ZN(
        \mult_x_9/n558 ) );
  NR2D0 U1879 ( .A1(n1742), .A2(n1529), .ZN(n1482) );
  OAI22D0 U1880 ( .A1(n1747), .A2(n1531), .B1(n1752), .B2(n1530), .ZN(n1481)
         );
  AOI211D0 U1881 ( .A1(n1745), .A2(n1534), .B(n1482), .C(n1481), .ZN(n1483) );
  MUX2ND0 U1882 ( .I0(R[17]), .I1(\mult_x_9/n556 ), .S(n1483), .ZN(
        \mult_x_9/n559 ) );
  NR2D0 U1883 ( .A1(n1747), .A2(n1529), .ZN(n1485) );
  OAI22D0 U1884 ( .A1(n1752), .A2(n1531), .B1(n1757), .B2(n1530), .ZN(n1484)
         );
  AOI211D0 U1885 ( .A1(n1750), .A2(n1534), .B(n1485), .C(n1484), .ZN(n1486) );
  MUX2ND0 U1886 ( .I0(R[17]), .I1(\mult_x_9/n556 ), .S(n1486), .ZN(
        \mult_x_9/n560 ) );
  NR2D0 U1887 ( .A1(n1752), .A2(n1529), .ZN(n1488) );
  OAI22D0 U1888 ( .A1(n1757), .A2(n1531), .B1(n1762), .B2(n1530), .ZN(n1487)
         );
  MUX2ND0 U1889 ( .I0(R[17]), .I1(\mult_x_9/n556 ), .S(n1489), .ZN(
        \mult_x_9/n561 ) );
  NR2D0 U1890 ( .A1(n1757), .A2(n1529), .ZN(n1491) );
  OAI22D0 U1891 ( .A1(n1762), .A2(n1531), .B1(n1767), .B2(n1530), .ZN(n1490)
         );
  AOI211D0 U1892 ( .A1(n1760), .A2(n1534), .B(n1491), .C(n1490), .ZN(n1492) );
  MUX2ND0 U1893 ( .I0(R[17]), .I1(\mult_x_9/n556 ), .S(n1492), .ZN(
        \mult_x_9/n562 ) );
  NR2D0 U1894 ( .A1(n1762), .A2(n1529), .ZN(n1494) );
  OAI22D0 U1895 ( .A1(n1767), .A2(n1531), .B1(n1772), .B2(n1530), .ZN(n1493)
         );
  AOI211D0 U1896 ( .A1(n1765), .A2(n1534), .B(n1494), .C(n1493), .ZN(n1495) );
  MUX2ND0 U1897 ( .I0(R[17]), .I1(\mult_x_9/n556 ), .S(n1495), .ZN(
        \mult_x_9/n563 ) );
  NR2D0 U1898 ( .A1(n1767), .A2(n1529), .ZN(n1497) );
  OAI22D0 U1899 ( .A1(n1772), .A2(n1531), .B1(n1777), .B2(n1530), .ZN(n1496)
         );
  AOI211D0 U1900 ( .A1(n1770), .A2(n1534), .B(n1497), .C(n1496), .ZN(n1498) );
  MUX2ND0 U1901 ( .I0(R[17]), .I1(\mult_x_9/n556 ), .S(n1498), .ZN(
        \mult_x_9/n564 ) );
  NR2D0 U1902 ( .A1(n1772), .A2(n1529), .ZN(n1500) );
  OAI22D0 U1903 ( .A1(n1777), .A2(n1531), .B1(n1782), .B2(n1530), .ZN(n1499)
         );
  AOI211D0 U1904 ( .A1(n1775), .A2(n1534), .B(n1500), .C(n1499), .ZN(n1501) );
  MUX2ND0 U1905 ( .I0(R[17]), .I1(\mult_x_9/n556 ), .S(n1501), .ZN(
        \mult_x_9/n565 ) );
  NR2D0 U1906 ( .A1(n1782), .A2(n1531), .ZN(n1503) );
  OAI22D0 U1907 ( .A1(n1777), .A2(n1529), .B1(n1787), .B2(n1530), .ZN(n1502)
         );
  AOI211D0 U1908 ( .A1(n1780), .A2(n1534), .B(n1503), .C(n1502), .ZN(n1504) );
  MUX2ND0 U1909 ( .I0(R[17]), .I1(\mult_x_9/n556 ), .S(n1504), .ZN(
        \mult_x_9/n566 ) );
  NR2D0 U1910 ( .A1(n1787), .A2(n1531), .ZN(n1506) );
  OAI22D0 U1911 ( .A1(n1782), .A2(n1529), .B1(n1792), .B2(n1530), .ZN(n1505)
         );
  AOI211D0 U1912 ( .A1(n1785), .A2(n1534), .B(n1506), .C(n1505), .ZN(n1507) );
  MUX2ND0 U1913 ( .I0(R[17]), .I1(\mult_x_9/n556 ), .S(n1507), .ZN(
        \mult_x_9/n567 ) );
  NR2D0 U1914 ( .A1(n1787), .A2(n1529), .ZN(n1509) );
  OAI22D0 U1915 ( .A1(n1792), .A2(n1531), .B1(n1797), .B2(n1530), .ZN(n1508)
         );
  AOI211D0 U1916 ( .A1(n1534), .A2(n1790), .B(n1509), .C(n1508), .ZN(n1510) );
  MUX2ND0 U1917 ( .I0(R[17]), .I1(\mult_x_9/n556 ), .S(n1510), .ZN(
        \mult_x_9/n568 ) );
  NR2D0 U1918 ( .A1(n1792), .A2(n1529), .ZN(n1512) );
  OAI22D0 U1919 ( .A1(n1797), .A2(n1531), .B1(n1802), .B2(n1530), .ZN(n1511)
         );
  AOI211D0 U1920 ( .A1(n1534), .A2(n1795), .B(n1512), .C(n1511), .ZN(n1513) );
  MUX2ND0 U1921 ( .I0(R[17]), .I1(\mult_x_9/n556 ), .S(n1513), .ZN(
        \mult_x_9/n569 ) );
  NR2D0 U1922 ( .A1(n1797), .A2(n1529), .ZN(n1515) );
  OAI22D0 U1923 ( .A1(n1802), .A2(n1531), .B1(n1807), .B2(n1530), .ZN(n1514)
         );
  AOI211D0 U1924 ( .A1(n1534), .A2(n1800), .B(n1515), .C(n1514), .ZN(n1516) );
  MUX2ND0 U1925 ( .I0(R[17]), .I1(\mult_x_9/n556 ), .S(n1516), .ZN(
        \mult_x_9/n570 ) );
  NR2D0 U1926 ( .A1(n1802), .A2(n1529), .ZN(n1518) );
  AOI211D0 U1927 ( .A1(n1534), .A2(n1805), .B(n1518), .C(n1517), .ZN(n1519) );
  MUX2ND0 U1928 ( .I0(R[17]), .I1(\mult_x_9/n556 ), .S(n1519), .ZN(
        \mult_x_9/n571 ) );
  NR2D0 U1929 ( .A1(n1807), .A2(n1529), .ZN(n1521) );
  OAI22D0 U1930 ( .A1(n1812), .A2(n1531), .B1(n1817), .B2(n1530), .ZN(n1520)
         );
  AOI211D0 U1931 ( .A1(n1534), .A2(n1810), .B(n1521), .C(n1520), .ZN(n1522) );
  MUX2ND0 U1932 ( .I0(R[17]), .I1(\mult_x_9/n556 ), .S(n1522), .ZN(
        \mult_x_9/n572 ) );
  NR2D0 U1933 ( .A1(n1812), .A2(n1529), .ZN(n1524) );
  OAI22D0 U1934 ( .A1(n1817), .A2(n1531), .B1(n1823), .B2(n1530), .ZN(n1523)
         );
  AOI211D0 U1935 ( .A1(n1534), .A2(n1815), .B(n1524), .C(n1523), .ZN(n1525) );
  MUX2ND0 U1936 ( .I0(R[17]), .I1(\mult_x_9/n556 ), .S(n1525), .ZN(
        \mult_x_9/n573 ) );
  NR2D0 U1937 ( .A1(n1817), .A2(n1529), .ZN(n1527) );
  OAI22D0 U1938 ( .A1(n1823), .A2(n1531), .B1(n1827), .B2(n1530), .ZN(n1526)
         );
  AOI211D0 U1939 ( .A1(n1534), .A2(n1820), .B(n1527), .C(n1526), .ZN(n1528) );
  MUX2ND0 U1940 ( .I0(R[17]), .I1(\mult_x_9/n556 ), .S(n1528), .ZN(
        \mult_x_9/n574 ) );
  OAI22D0 U1941 ( .A1(n1827), .A2(n1531), .B1(n1825), .B2(n1530), .ZN(n1532)
         );
  AOI211D0 U1942 ( .A1(n1534), .A2(n1831), .B(n1533), .C(n1532), .ZN(n1535) );
  MUX2ND0 U1943 ( .I0(R[17]), .I1(\mult_x_9/n556 ), .S(n1535), .ZN(
        \mult_x_9/n575 ) );
  OAI22D0 U1944 ( .A1(n1742), .A2(n1597), .B1(n1537), .B2(n1737), .ZN(n1536)
         );
  MUX2ND0 U1945 ( .I0(n1603), .I1(R[14]), .S(n1536), .ZN(\mult_x_9/n583 ) );
  OAI222D0 U1946 ( .A1(n1739), .A2(n1537), .B1(n1596), .B2(n1742), .C1(n1597), 
        .C2(n1747), .ZN(n1538) );
  MUX2ND0 U1947 ( .I0(n1603), .I1(R[14]), .S(n1538), .ZN(\mult_x_9/n584 ) );
  NR2D0 U1948 ( .A1(n1747), .A2(n1596), .ZN(n1540) );
  OAI22D0 U1949 ( .A1(n1742), .A2(n1598), .B1(n1752), .B2(n1597), .ZN(n1539)
         );
  AOI211D0 U1950 ( .A1(n1745), .A2(n1601), .B(n1540), .C(n1539), .ZN(n1541) );
  MUX2ND0 U1951 ( .I0(R[14]), .I1(n1603), .S(n1541), .ZN(\mult_x_9/n585 ) );
  NR2D0 U1952 ( .A1(n1752), .A2(n1596), .ZN(n1543) );
  AOI211D0 U1953 ( .A1(n1750), .A2(n1601), .B(n1543), .C(n1542), .ZN(n1544) );
  MUX2ND0 U1954 ( .I0(R[14]), .I1(n1603), .S(n1544), .ZN(\mult_x_9/n586 ) );
  NR2D0 U1955 ( .A1(n1757), .A2(n1596), .ZN(n1546) );
  OAI22D0 U1956 ( .A1(n1752), .A2(n1598), .B1(n1762), .B2(n1597), .ZN(n1545)
         );
  AOI211D0 U1957 ( .A1(n1755), .A2(n1601), .B(n1546), .C(n1545), .ZN(n1547) );
  MUX2ND0 U1958 ( .I0(R[14]), .I1(n1603), .S(n1547), .ZN(\mult_x_9/n587 ) );
  NR2D0 U1959 ( .A1(n1762), .A2(n1596), .ZN(n1549) );
  OAI22D0 U1960 ( .A1(n1757), .A2(n1598), .B1(n1767), .B2(n1597), .ZN(n1548)
         );
  AOI211D0 U1961 ( .A1(n1760), .A2(n1601), .B(n1549), .C(n1548), .ZN(n1550) );
  MUX2ND0 U1962 ( .I0(R[14]), .I1(n1603), .S(n1550), .ZN(\mult_x_9/n588 ) );
  OAI22D0 U1963 ( .A1(n1762), .A2(n1598), .B1(n1772), .B2(n1597), .ZN(n1551)
         );
  AOI211D0 U1964 ( .A1(n1765), .A2(n1601), .B(n1552), .C(n1551), .ZN(n1553) );
  MUX2ND0 U1965 ( .I0(R[14]), .I1(n1603), .S(n1553), .ZN(\mult_x_9/n589 ) );
  NR2D0 U1966 ( .A1(n1772), .A2(n1596), .ZN(n1555) );
  OAI22D0 U1967 ( .A1(n1767), .A2(n1598), .B1(n1777), .B2(n1597), .ZN(n1554)
         );
  AOI211D0 U1968 ( .A1(n1770), .A2(n1601), .B(n1555), .C(n1554), .ZN(n1556) );
  MUX2ND0 U1969 ( .I0(R[14]), .I1(n1603), .S(n1556), .ZN(\mult_x_9/n590 ) );
  NR2D0 U1970 ( .A1(n1777), .A2(n1596), .ZN(n1558) );
  OAI22D0 U1971 ( .A1(n1772), .A2(n1598), .B1(n1782), .B2(n1597), .ZN(n1557)
         );
  AOI211D0 U1972 ( .A1(n1775), .A2(n1601), .B(n1558), .C(n1557), .ZN(n1559) );
  MUX2ND0 U1973 ( .I0(R[14]), .I1(n1603), .S(n1559), .ZN(\mult_x_9/n591 ) );
  NR2D0 U1974 ( .A1(n1787), .A2(n1597), .ZN(n1561) );
  OAI22D0 U1975 ( .A1(n1777), .A2(n1598), .B1(n1782), .B2(n1596), .ZN(n1560)
         );
  AOI211D0 U1976 ( .A1(n1780), .A2(n1601), .B(n1561), .C(n1560), .ZN(n1562) );
  MUX2ND0 U1977 ( .I0(R[14]), .I1(n1603), .S(n1562), .ZN(\mult_x_9/n592 ) );
  NR2D0 U1978 ( .A1(n1792), .A2(n1597), .ZN(n1564) );
  OAI22D0 U1979 ( .A1(n1782), .A2(n1598), .B1(n1787), .B2(n1596), .ZN(n1563)
         );
  AOI211D0 U1980 ( .A1(n1785), .A2(n1601), .B(n1564), .C(n1563), .ZN(n1565) );
  MUX2ND0 U1981 ( .I0(R[14]), .I1(n1603), .S(n1565), .ZN(\mult_x_9/n593 ) );
  NR2D0 U1982 ( .A1(n1792), .A2(n1596), .ZN(n1567) );
  OAI22D0 U1983 ( .A1(n1787), .A2(n1598), .B1(n1797), .B2(n1597), .ZN(n1566)
         );
  AOI211D0 U1984 ( .A1(n1601), .A2(n1790), .B(n1567), .C(n1566), .ZN(n1568) );
  MUX2ND0 U1985 ( .I0(R[14]), .I1(n1603), .S(n1568), .ZN(\mult_x_9/n594 ) );
  OAI22D0 U1986 ( .A1(n1792), .A2(n1598), .B1(n1802), .B2(n1597), .ZN(n1569)
         );
  AOI211D0 U1987 ( .A1(n1601), .A2(n1795), .B(n1570), .C(n1569), .ZN(n1571) );
  MUX2ND0 U1988 ( .I0(R[14]), .I1(n1603), .S(n1571), .ZN(\mult_x_9/n595 ) );
  NR2D0 U1989 ( .A1(n1802), .A2(n1596), .ZN(n1573) );
  OAI22D0 U1990 ( .A1(n1797), .A2(n1598), .B1(n1807), .B2(n1597), .ZN(n1572)
         );
  AOI211D0 U1991 ( .A1(n1601), .A2(n1800), .B(n1573), .C(n1572), .ZN(n1574) );
  MUX2ND0 U1992 ( .I0(R[14]), .I1(n1603), .S(n1574), .ZN(\mult_x_9/n596 ) );
  NR2D0 U1993 ( .A1(n1807), .A2(n1596), .ZN(n1576) );
  OAI22D0 U1994 ( .A1(n1802), .A2(n1598), .B1(n1812), .B2(n1597), .ZN(n1575)
         );
  AOI211D0 U1995 ( .A1(n1601), .A2(n1805), .B(n1576), .C(n1575), .ZN(n1577) );
  MUX2ND0 U1996 ( .I0(R[14]), .I1(n1603), .S(n1577), .ZN(\mult_x_9/n597 ) );
  NR2D0 U1997 ( .A1(n1812), .A2(n1596), .ZN(n1579) );
  OAI22D0 U1998 ( .A1(n1807), .A2(n1598), .B1(n1817), .B2(n1597), .ZN(n1578)
         );
  AOI211D0 U1999 ( .A1(n1601), .A2(n1810), .B(n1579), .C(n1578), .ZN(n1580) );
  MUX2ND0 U2000 ( .I0(R[14]), .I1(n1603), .S(n1580), .ZN(\mult_x_9/n598 ) );
  NR2D0 U2001 ( .A1(n1817), .A2(n1596), .ZN(n1582) );
  OAI22D0 U2002 ( .A1(n1812), .A2(n1598), .B1(n1823), .B2(n1597), .ZN(n1581)
         );
  AOI211D0 U2003 ( .A1(n1601), .A2(n1815), .B(n1582), .C(n1581), .ZN(n1583) );
  MUX2ND0 U2004 ( .I0(R[14]), .I1(n1603), .S(n1583), .ZN(\mult_x_9/n599 ) );
  OAI22D0 U2005 ( .A1(n1817), .A2(n1598), .B1(n1827), .B2(n1597), .ZN(n1584)
         );
  AOI211D0 U2006 ( .A1(n1601), .A2(n1820), .B(n1585), .C(n1584), .ZN(n1586) );
  MUX2ND0 U2007 ( .I0(R[14]), .I1(n1603), .S(n1586), .ZN(\mult_x_9/n600 ) );
  NR2D0 U2008 ( .A1(n1827), .A2(n1596), .ZN(n1588) );
  OAI22D0 U2009 ( .A1(n1823), .A2(n1598), .B1(n1825), .B2(n1597), .ZN(n1587)
         );
  AOI211D0 U2010 ( .A1(n1601), .A2(n1831), .B(n1588), .C(n1587), .ZN(n1589) );
  MUX2ND0 U2011 ( .I0(R[14]), .I1(n1603), .S(n1589), .ZN(\mult_x_9/n601 ) );
  NR2D0 U2012 ( .A1(n1825), .A2(n1596), .ZN(n1591) );
  OAI22D0 U2013 ( .A1(n1827), .A2(n1598), .B1(n1730), .B2(n1597), .ZN(n1590)
         );
  AOI211D0 U2014 ( .A1(n1601), .A2(n1719), .B(n1591), .C(n1590), .ZN(n1592) );
  MUX2ND0 U2015 ( .I0(R[14]), .I1(n1603), .S(n1592), .ZN(\mult_x_9/n602 ) );
  NR2D0 U2016 ( .A1(n1730), .A2(n1596), .ZN(n1594) );
  OAI22D0 U2017 ( .A1(n1825), .A2(n1598), .B1(n1726), .B2(n1597), .ZN(n1593)
         );
  AOI211D0 U2018 ( .A1(n1601), .A2(n1723), .B(n1594), .C(n1593), .ZN(n1595) );
  MUX2ND0 U2019 ( .I0(R[14]), .I1(n1603), .S(n1595), .ZN(\mult_x_9/n603 ) );
  NR2D0 U2020 ( .A1(n1726), .A2(n1596), .ZN(n1600) );
  OAI22D0 U2021 ( .A1(n1730), .A2(n1598), .B1(n1728), .B2(n1597), .ZN(n1599)
         );
  AOI211D0 U2022 ( .A1(n1601), .A2(n1733), .B(n1600), .C(n1599), .ZN(n1602) );
  MUX2ND0 U2023 ( .I0(R[14]), .I1(n1603), .S(n1602), .ZN(\mult_x_9/n604 ) );
  OAI22D0 U2024 ( .A1(n1742), .A2(n1656), .B1(n1605), .B2(n1737), .ZN(n1604)
         );
  MUX2ND0 U2025 ( .I0(\mult_x_9/n608 ), .I1(R[11]), .S(n1604), .ZN(
        \mult_x_9/n609 ) );
  OAI222D0 U2026 ( .A1(n1656), .A2(n1747), .B1(n1657), .B2(n1742), .C1(n1605), 
        .C2(n1739), .ZN(n1606) );
  MUX2ND0 U2027 ( .I0(\mult_x_9/n608 ), .I1(R[11]), .S(n1606), .ZN(
        \mult_x_9/n610 ) );
  NR2D0 U2028 ( .A1(n1742), .A2(n1655), .ZN(n1608) );
  OAI22D0 U2029 ( .A1(n1747), .A2(n1657), .B1(n1752), .B2(n1656), .ZN(n1607)
         );
  AOI211D0 U2030 ( .A1(n1745), .A2(n1660), .B(n1608), .C(n1607), .ZN(n1609) );
  MUX2ND0 U2031 ( .I0(R[11]), .I1(\mult_x_9/n608 ), .S(n1609), .ZN(
        \mult_x_9/n611 ) );
  NR2D0 U2032 ( .A1(n1747), .A2(n1655), .ZN(n1611) );
  OAI22D0 U2033 ( .A1(n1752), .A2(n1657), .B1(n1757), .B2(n1656), .ZN(n1610)
         );
  AOI211D0 U2034 ( .A1(n1750), .A2(n1660), .B(n1611), .C(n1610), .ZN(n1612) );
  MUX2ND0 U2035 ( .I0(R[11]), .I1(\mult_x_9/n608 ), .S(n1612), .ZN(
        \mult_x_9/n612 ) );
  NR2D0 U2036 ( .A1(n1752), .A2(n1655), .ZN(n1614) );
  AOI211D0 U2037 ( .A1(n1755), .A2(n1660), .B(n1614), .C(n1613), .ZN(n1615) );
  MUX2ND0 U2038 ( .I0(R[11]), .I1(\mult_x_9/n608 ), .S(n1615), .ZN(
        \mult_x_9/n613 ) );
  NR2D0 U2039 ( .A1(n1757), .A2(n1655), .ZN(n1617) );
  OAI22D0 U2040 ( .A1(n1762), .A2(n1657), .B1(n1767), .B2(n1656), .ZN(n1616)
         );
  AOI211D0 U2041 ( .A1(n1760), .A2(n1660), .B(n1617), .C(n1616), .ZN(n1618) );
  MUX2ND0 U2042 ( .I0(R[11]), .I1(\mult_x_9/n608 ), .S(n1618), .ZN(
        \mult_x_9/n614 ) );
  NR2D0 U2043 ( .A1(n1762), .A2(n1655), .ZN(n1620) );
  OAI22D0 U2044 ( .A1(n1767), .A2(n1657), .B1(n1772), .B2(n1656), .ZN(n1619)
         );
  AOI211D0 U2045 ( .A1(n1765), .A2(n1660), .B(n1620), .C(n1619), .ZN(n1621) );
  MUX2ND0 U2046 ( .I0(R[11]), .I1(\mult_x_9/n608 ), .S(n1621), .ZN(
        \mult_x_9/n615 ) );
  NR2D0 U2047 ( .A1(n1767), .A2(n1655), .ZN(n1623) );
  MUX2ND0 U2048 ( .I0(R[11]), .I1(\mult_x_9/n608 ), .S(n1624), .ZN(
        \mult_x_9/n616 ) );
  NR2D0 U2049 ( .A1(n1772), .A2(n1655), .ZN(n1626) );
  OAI22D0 U2050 ( .A1(n1777), .A2(n1657), .B1(n1782), .B2(n1656), .ZN(n1625)
         );
  AOI211D0 U2051 ( .A1(n1775), .A2(n1660), .B(n1626), .C(n1625), .ZN(n1627) );
  MUX2ND0 U2052 ( .I0(R[11]), .I1(\mult_x_9/n608 ), .S(n1627), .ZN(
        \mult_x_9/n617 ) );
  NR2D0 U2053 ( .A1(n1782), .A2(n1657), .ZN(n1629) );
  OAI22D0 U2054 ( .A1(n1777), .A2(n1655), .B1(n1787), .B2(n1656), .ZN(n1628)
         );
  AOI211D0 U2055 ( .A1(n1780), .A2(n1660), .B(n1629), .C(n1628), .ZN(n1630) );
  MUX2ND0 U2056 ( .I0(R[11]), .I1(\mult_x_9/n608 ), .S(n1630), .ZN(
        \mult_x_9/n618 ) );
  NR2D0 U2057 ( .A1(n1787), .A2(n1657), .ZN(n1632) );
  OAI22D0 U2058 ( .A1(n1782), .A2(n1655), .B1(n1792), .B2(n1656), .ZN(n1631)
         );
  MUX2ND0 U2059 ( .I0(R[11]), .I1(\mult_x_9/n608 ), .S(n1633), .ZN(
        \mult_x_9/n619 ) );
  NR2D0 U2060 ( .A1(n1787), .A2(n1655), .ZN(n1635) );
  OAI22D0 U2061 ( .A1(n1792), .A2(n1657), .B1(n1797), .B2(n1656), .ZN(n1634)
         );
  AOI211D0 U2062 ( .A1(n1660), .A2(n1790), .B(n1635), .C(n1634), .ZN(n1636) );
  MUX2ND0 U2063 ( .I0(R[11]), .I1(\mult_x_9/n608 ), .S(n1636), .ZN(
        \mult_x_9/n620 ) );
  NR2D0 U2064 ( .A1(n1792), .A2(n1655), .ZN(n1638) );
  OAI22D0 U2065 ( .A1(n1797), .A2(n1657), .B1(n1802), .B2(n1656), .ZN(n1637)
         );
  AOI211D0 U2066 ( .A1(n1660), .A2(n1795), .B(n1638), .C(n1637), .ZN(n1639) );
  MUX2ND0 U2067 ( .I0(R[11]), .I1(\mult_x_9/n608 ), .S(n1639), .ZN(
        \mult_x_9/n621 ) );
  NR2D0 U2068 ( .A1(n1797), .A2(n1655), .ZN(n1641) );
  OAI22D0 U2069 ( .A1(n1802), .A2(n1657), .B1(n1807), .B2(n1656), .ZN(n1640)
         );
  AOI211D0 U2070 ( .A1(n1660), .A2(n1800), .B(n1641), .C(n1640), .ZN(n1642) );
  MUX2ND0 U2071 ( .I0(R[11]), .I1(\mult_x_9/n608 ), .S(n1642), .ZN(
        \mult_x_9/n622 ) );
  NR2D0 U2072 ( .A1(n1802), .A2(n1655), .ZN(n1644) );
  OAI22D0 U2073 ( .A1(n1807), .A2(n1657), .B1(n1812), .B2(n1656), .ZN(n1643)
         );
  AOI211D0 U2074 ( .A1(n1660), .A2(n1805), .B(n1644), .C(n1643), .ZN(n1645) );
  MUX2ND0 U2075 ( .I0(R[11]), .I1(\mult_x_9/n608 ), .S(n1645), .ZN(
        \mult_x_9/n623 ) );
  NR2D0 U2076 ( .A1(n1807), .A2(n1655), .ZN(n1647) );
  OAI22D0 U2077 ( .A1(n1812), .A2(n1657), .B1(n1817), .B2(n1656), .ZN(n1646)
         );
  AOI211D0 U2078 ( .A1(n1660), .A2(n1810), .B(n1647), .C(n1646), .ZN(n1648) );
  MUX2ND0 U2079 ( .I0(R[11]), .I1(\mult_x_9/n608 ), .S(n1648), .ZN(
        \mult_x_9/n624 ) );
  OAI22D0 U2080 ( .A1(n1817), .A2(n1657), .B1(n1823), .B2(n1656), .ZN(n1649)
         );
  AOI211D0 U2081 ( .A1(n1660), .A2(n1815), .B(n1650), .C(n1649), .ZN(n1651) );
  MUX2ND0 U2082 ( .I0(R[11]), .I1(\mult_x_9/n608 ), .S(n1651), .ZN(
        \mult_x_9/n625 ) );
  NR2D0 U2083 ( .A1(n1817), .A2(n1655), .ZN(n1653) );
  OAI22D0 U2084 ( .A1(n1823), .A2(n1657), .B1(n1827), .B2(n1656), .ZN(n1652)
         );
  AOI211D0 U2085 ( .A1(n1660), .A2(n1820), .B(n1653), .C(n1652), .ZN(n1654) );
  MUX2ND0 U2086 ( .I0(R[11]), .I1(\mult_x_9/n608 ), .S(n1654), .ZN(
        \mult_x_9/n626 ) );
  NR2D0 U2087 ( .A1(n1823), .A2(n1655), .ZN(n1659) );
  OAI22D0 U2088 ( .A1(n1827), .A2(n1657), .B1(n1825), .B2(n1656), .ZN(n1658)
         );
  AOI211D0 U2089 ( .A1(n1660), .A2(n1831), .B(n1659), .C(n1658), .ZN(n1661) );
  MUX2ND0 U2090 ( .I0(R[11]), .I1(\mult_x_9/n608 ), .S(n1661), .ZN(
        \mult_x_9/n627 ) );
  INVD0 U2091 ( .I(n1662), .ZN(n1727) );
  OAI22D0 U2092 ( .A1(n1742), .A2(n1727), .B1(n1664), .B2(n1737), .ZN(n1663)
         );
  MUX2ND0 U2093 ( .I0(n1736), .I1(R[8]), .S(n1663), .ZN(\mult_x_9/n635 ) );
  OAI222D0 U2094 ( .A1(n1727), .A2(n1747), .B1(n1725), .B2(n1742), .C1(n1664), 
        .C2(n1739), .ZN(n1665) );
  MUX2ND0 U2095 ( .I0(n1736), .I1(R[8]), .S(n1665), .ZN(\mult_x_9/n636 ) );
  NR2D0 U2096 ( .A1(n1747), .A2(n1725), .ZN(n1667) );
  OAI22D0 U2097 ( .A1(n1742), .A2(n1729), .B1(n1752), .B2(n1727), .ZN(n1666)
         );
  AOI211D0 U2098 ( .A1(n1745), .A2(n1734), .B(n1667), .C(n1666), .ZN(n1668) );
  MUX2ND0 U2099 ( .I0(R[8]), .I1(n1736), .S(n1668), .ZN(\mult_x_9/n637 ) );
  NR2D0 U2100 ( .A1(n1752), .A2(n1725), .ZN(n1670) );
  OAI22D0 U2101 ( .A1(n1747), .A2(n1729), .B1(n1757), .B2(n1727), .ZN(n1669)
         );
  AOI211D0 U2102 ( .A1(n1750), .A2(n1734), .B(n1670), .C(n1669), .ZN(n1671) );
  MUX2ND0 U2103 ( .I0(R[8]), .I1(n1736), .S(n1671), .ZN(\mult_x_9/n638 ) );
  NR2D0 U2104 ( .A1(n1757), .A2(n1725), .ZN(n1673) );
  OAI22D0 U2105 ( .A1(n1752), .A2(n1729), .B1(n1762), .B2(n1727), .ZN(n1672)
         );
  AOI211D0 U2106 ( .A1(n1755), .A2(n1734), .B(n1673), .C(n1672), .ZN(n1674) );
  MUX2ND0 U2107 ( .I0(R[8]), .I1(n1736), .S(n1674), .ZN(\mult_x_9/n639 ) );
  NR2D0 U2108 ( .A1(n1762), .A2(n1725), .ZN(n1676) );
  OAI22D0 U2109 ( .A1(n1757), .A2(n1729), .B1(n1767), .B2(n1727), .ZN(n1675)
         );
  AOI211D0 U2110 ( .A1(n1760), .A2(n1734), .B(n1676), .C(n1675), .ZN(n1677) );
  MUX2ND0 U2111 ( .I0(R[8]), .I1(n1736), .S(n1677), .ZN(\mult_x_9/n640 ) );
  NR2D0 U2112 ( .A1(n1767), .A2(n1725), .ZN(n1679) );
  OAI22D0 U2113 ( .A1(n1762), .A2(n1729), .B1(n1772), .B2(n1727), .ZN(n1678)
         );
  AOI211D0 U2114 ( .A1(n1765), .A2(n1734), .B(n1679), .C(n1678), .ZN(n1680) );
  MUX2ND0 U2115 ( .I0(R[8]), .I1(n1736), .S(n1680), .ZN(\mult_x_9/n641 ) );
  NR2D0 U2116 ( .A1(n1772), .A2(n1725), .ZN(n1682) );
  OAI22D0 U2117 ( .A1(n1767), .A2(n1729), .B1(n1777), .B2(n1727), .ZN(n1681)
         );
  AOI211D0 U2118 ( .A1(n1770), .A2(n1734), .B(n1682), .C(n1681), .ZN(n1683) );
  MUX2ND0 U2119 ( .I0(R[8]), .I1(n1736), .S(n1683), .ZN(\mult_x_9/n642 ) );
  NR2D0 U2120 ( .A1(n1777), .A2(n1725), .ZN(n1685) );
  OAI22D0 U2121 ( .A1(n1772), .A2(n1729), .B1(n1782), .B2(n1727), .ZN(n1684)
         );
  AOI211D0 U2122 ( .A1(n1775), .A2(n1734), .B(n1685), .C(n1684), .ZN(n1686) );
  MUX2ND0 U2123 ( .I0(R[8]), .I1(n1736), .S(n1686), .ZN(\mult_x_9/n643 ) );
  NR2D0 U2124 ( .A1(n1787), .A2(n1727), .ZN(n1688) );
  OAI22D0 U2125 ( .A1(n1777), .A2(n1729), .B1(n1782), .B2(n1725), .ZN(n1687)
         );
  AOI211D0 U2126 ( .A1(n1780), .A2(n1734), .B(n1688), .C(n1687), .ZN(n1689) );
  MUX2ND0 U2127 ( .I0(R[8]), .I1(n1736), .S(n1689), .ZN(\mult_x_9/n644 ) );
  NR2D0 U2128 ( .A1(n1792), .A2(n1727), .ZN(n1691) );
  OAI22D0 U2129 ( .A1(n1782), .A2(n1729), .B1(n1787), .B2(n1725), .ZN(n1690)
         );
  AOI211D0 U2130 ( .A1(n1785), .A2(n1734), .B(n1691), .C(n1690), .ZN(n1692) );
  MUX2ND0 U2131 ( .I0(R[8]), .I1(n1736), .S(n1692), .ZN(\mult_x_9/n645 ) );
  NR2D0 U2132 ( .A1(n1792), .A2(n1725), .ZN(n1694) );
  OAI22D0 U2133 ( .A1(n1787), .A2(n1729), .B1(n1797), .B2(n1727), .ZN(n1693)
         );
  AOI211D0 U2134 ( .A1(n1734), .A2(n1790), .B(n1694), .C(n1693), .ZN(n1695) );
  MUX2ND0 U2135 ( .I0(R[8]), .I1(n1736), .S(n1695), .ZN(\mult_x_9/n646 ) );
  NR2D0 U2136 ( .A1(n1797), .A2(n1725), .ZN(n1697) );
  AOI211D0 U2137 ( .A1(n1734), .A2(n1795), .B(n1697), .C(n1696), .ZN(n1698) );
  MUX2ND0 U2138 ( .I0(R[8]), .I1(n1736), .S(n1698), .ZN(\mult_x_9/n647 ) );
  NR2D0 U2139 ( .A1(n1802), .A2(n1725), .ZN(n1700) );
  OAI22D0 U2140 ( .A1(n1797), .A2(n1729), .B1(n1807), .B2(n1727), .ZN(n1699)
         );
  AOI211D0 U2141 ( .A1(n1734), .A2(n1800), .B(n1700), .C(n1699), .ZN(n1701) );
  MUX2ND0 U2142 ( .I0(R[8]), .I1(n1736), .S(n1701), .ZN(\mult_x_9/n648 ) );
  OAI22D0 U2143 ( .A1(n1802), .A2(n1729), .B1(n1812), .B2(n1727), .ZN(n1702)
         );
  AOI211D0 U2144 ( .A1(n1734), .A2(n1805), .B(n1703), .C(n1702), .ZN(n1704) );
  MUX2ND0 U2145 ( .I0(R[8]), .I1(n1736), .S(n1704), .ZN(\mult_x_9/n649 ) );
  NR2D0 U2146 ( .A1(n1812), .A2(n1725), .ZN(n1706) );
  OAI22D0 U2147 ( .A1(n1807), .A2(n1729), .B1(n1817), .B2(n1727), .ZN(n1705)
         );
  AOI211D0 U2148 ( .A1(n1734), .A2(n1810), .B(n1706), .C(n1705), .ZN(n1707) );
  MUX2ND0 U2149 ( .I0(R[8]), .I1(n1736), .S(n1707), .ZN(\mult_x_9/n650 ) );
  NR2D0 U2150 ( .A1(n1817), .A2(n1725), .ZN(n1709) );
  OAI22D0 U2151 ( .A1(n1812), .A2(n1729), .B1(n1823), .B2(n1727), .ZN(n1708)
         );
  AOI211D0 U2152 ( .A1(n1734), .A2(n1815), .B(n1709), .C(n1708), .ZN(n1710) );
  MUX2ND0 U2153 ( .I0(R[8]), .I1(n1736), .S(n1710), .ZN(\mult_x_9/n651 ) );
  NR2D0 U2154 ( .A1(n1823), .A2(n1725), .ZN(n1712) );
  AOI211D0 U2155 ( .A1(n1734), .A2(n1820), .B(n1712), .C(n1711), .ZN(n1713) );
  MUX2ND0 U2156 ( .I0(R[8]), .I1(n1736), .S(n1713), .ZN(\mult_x_9/n652 ) );
  NR2D0 U2157 ( .A1(n1827), .A2(n1725), .ZN(n1715) );
  AOI211D0 U2158 ( .A1(n1734), .A2(n1831), .B(n1715), .C(n1714), .ZN(n1716) );
  MUX2ND0 U2159 ( .I0(R[8]), .I1(n1736), .S(n1716), .ZN(\mult_x_9/n653 ) );
  NR2D0 U2160 ( .A1(n1825), .A2(n1725), .ZN(n1718) );
  OAI22D0 U2161 ( .A1(n1827), .A2(n1729), .B1(n1730), .B2(n1727), .ZN(n1717)
         );
  AOI211D0 U2162 ( .A1(n1734), .A2(n1719), .B(n1718), .C(n1717), .ZN(n1720) );
  MUX2ND0 U2163 ( .I0(R[8]), .I1(n1736), .S(n1720), .ZN(\mult_x_9/n654 ) );
  NR2D0 U2164 ( .A1(n1730), .A2(n1725), .ZN(n1722) );
  OAI22D0 U2165 ( .A1(n1825), .A2(n1729), .B1(n1726), .B2(n1727), .ZN(n1721)
         );
  AOI211D0 U2166 ( .A1(n1734), .A2(n1723), .B(n1722), .C(n1721), .ZN(n1724) );
  MUX2ND0 U2167 ( .I0(R[8]), .I1(n1736), .S(n1724), .ZN(\mult_x_9/n655 ) );
  NR2D0 U2168 ( .A1(n1726), .A2(n1725), .ZN(n1732) );
  OAI22D0 U2169 ( .A1(n1730), .A2(n1729), .B1(n1728), .B2(n1727), .ZN(n1731)
         );
  AOI211D0 U2170 ( .A1(n1734), .A2(n1733), .B(n1732), .C(n1731), .ZN(n1735) );
  MUX2ND0 U2171 ( .I0(R[8]), .I1(n1736), .S(n1735), .ZN(\mult_x_9/n656 ) );
  OAI22D0 U2172 ( .A1(n1742), .A2(n1824), .B1(n1740), .B2(n1737), .ZN(n1738)
         );
  MUX2ND0 U2173 ( .I0(\mult_x_9/n660 ), .I1(R[5]), .S(n1738), .ZN(
        \mult_x_9/n661 ) );
  OAI222D0 U2174 ( .A1(n1824), .A2(n1747), .B1(n1826), .B2(n1742), .C1(n1740), 
        .C2(n1739), .ZN(n1741) );
  MUX2ND0 U2175 ( .I0(\mult_x_9/n660 ), .I1(R[5]), .S(n1741), .ZN(
        \mult_x_9/n662 ) );
  NR2D0 U2176 ( .A1(n1742), .A2(n1822), .ZN(n1744) );
  OAI22D0 U2177 ( .A1(n1747), .A2(n1826), .B1(n1752), .B2(n1824), .ZN(n1743)
         );
  AOI211D0 U2178 ( .A1(n1745), .A2(n1830), .B(n1744), .C(n1743), .ZN(n1746) );
  MUX2ND0 U2179 ( .I0(R[5]), .I1(\mult_x_9/n660 ), .S(n1746), .ZN(
        \mult_x_9/n663 ) );
  NR2D0 U2180 ( .A1(n1747), .A2(n1822), .ZN(n1749) );
  OAI22D0 U2181 ( .A1(n1752), .A2(n1826), .B1(n1757), .B2(n1824), .ZN(n1748)
         );
  MUX2ND0 U2182 ( .I0(R[5]), .I1(\mult_x_9/n660 ), .S(n1751), .ZN(
        \mult_x_9/n664 ) );
  NR2D0 U2183 ( .A1(n1752), .A2(n1822), .ZN(n1754) );
  OAI22D0 U2184 ( .A1(n1757), .A2(n1826), .B1(n1762), .B2(n1824), .ZN(n1753)
         );
  AOI211D0 U2185 ( .A1(n1755), .A2(n1830), .B(n1754), .C(n1753), .ZN(n1756) );
  MUX2ND0 U2186 ( .I0(R[5]), .I1(\mult_x_9/n660 ), .S(n1756), .ZN(
        \mult_x_9/n665 ) );
  NR2D0 U2187 ( .A1(n1757), .A2(n1822), .ZN(n1759) );
  OAI22D0 U2188 ( .A1(n1762), .A2(n1826), .B1(n1767), .B2(n1824), .ZN(n1758)
         );
  AOI211D0 U2189 ( .A1(n1760), .A2(n1830), .B(n1759), .C(n1758), .ZN(n1761) );
  MUX2ND0 U2190 ( .I0(R[5]), .I1(\mult_x_9/n660 ), .S(n1761), .ZN(
        \mult_x_9/n666 ) );
  NR2D0 U2191 ( .A1(n1762), .A2(n1822), .ZN(n1764) );
  OAI22D0 U2192 ( .A1(n1767), .A2(n1826), .B1(n1772), .B2(n1824), .ZN(n1763)
         );
  AOI211D0 U2193 ( .A1(n1765), .A2(n1830), .B(n1764), .C(n1763), .ZN(n1766) );
  MUX2ND0 U2194 ( .I0(R[5]), .I1(\mult_x_9/n660 ), .S(n1766), .ZN(
        \mult_x_9/n667 ) );
  OAI22D0 U2195 ( .A1(n1772), .A2(n1826), .B1(n1777), .B2(n1824), .ZN(n1768)
         );
  AOI211D0 U2196 ( .A1(n1770), .A2(n1830), .B(n1769), .C(n1768), .ZN(n1771) );
  MUX2ND0 U2197 ( .I0(R[5]), .I1(\mult_x_9/n660 ), .S(n1771), .ZN(
        \mult_x_9/n668 ) );
  NR2D0 U2198 ( .A1(n1772), .A2(n1822), .ZN(n1774) );
  OAI22D0 U2199 ( .A1(n1777), .A2(n1826), .B1(n1782), .B2(n1824), .ZN(n1773)
         );
  AOI211D0 U2200 ( .A1(n1775), .A2(n1830), .B(n1774), .C(n1773), .ZN(n1776) );
  MUX2ND0 U2201 ( .I0(R[5]), .I1(\mult_x_9/n660 ), .S(n1776), .ZN(
        \mult_x_9/n669 ) );
  NR2D0 U2202 ( .A1(n1782), .A2(n1826), .ZN(n1779) );
  OAI22D0 U2203 ( .A1(n1777), .A2(n1822), .B1(n1787), .B2(n1824), .ZN(n1778)
         );
  AOI211D0 U2204 ( .A1(n1780), .A2(n1830), .B(n1779), .C(n1778), .ZN(n1781) );
  MUX2ND0 U2205 ( .I0(R[5]), .I1(\mult_x_9/n660 ), .S(n1781), .ZN(
        \mult_x_9/n670 ) );
  NR2D0 U2206 ( .A1(n1787), .A2(n1826), .ZN(n1784) );
  OAI22D0 U2207 ( .A1(n1782), .A2(n1822), .B1(n1792), .B2(n1824), .ZN(n1783)
         );
  AOI211D0 U2208 ( .A1(n1785), .A2(n1830), .B(n1784), .C(n1783), .ZN(n1786) );
  MUX2ND0 U2209 ( .I0(R[5]), .I1(\mult_x_9/n660 ), .S(n1786), .ZN(
        \mult_x_9/n671 ) );
  NR2D0 U2210 ( .A1(n1787), .A2(n1822), .ZN(n1789) );
  OAI22D0 U2211 ( .A1(n1792), .A2(n1826), .B1(n1797), .B2(n1824), .ZN(n1788)
         );
  AOI211D0 U2212 ( .A1(n1790), .A2(n1830), .B(n1789), .C(n1788), .ZN(n1791) );
  MUX2ND0 U2213 ( .I0(R[5]), .I1(\mult_x_9/n660 ), .S(n1791), .ZN(
        \mult_x_9/n672 ) );
  NR2D0 U2214 ( .A1(n1792), .A2(n1822), .ZN(n1794) );
  OAI22D0 U2215 ( .A1(n1797), .A2(n1826), .B1(n1802), .B2(n1824), .ZN(n1793)
         );
  AOI211D0 U2216 ( .A1(n1795), .A2(n1830), .B(n1794), .C(n1793), .ZN(n1796) );
  MUX2ND0 U2217 ( .I0(R[5]), .I1(\mult_x_9/n660 ), .S(n1796), .ZN(
        \mult_x_9/n673 ) );
  NR2D0 U2218 ( .A1(n1797), .A2(n1822), .ZN(n1799) );
  OAI22D0 U2219 ( .A1(n1802), .A2(n1826), .B1(n1807), .B2(n1824), .ZN(n1798)
         );
  AOI211D0 U2220 ( .A1(n1800), .A2(n1830), .B(n1799), .C(n1798), .ZN(n1801) );
  MUX2ND0 U2221 ( .I0(R[5]), .I1(\mult_x_9/n660 ), .S(n1801), .ZN(
        \mult_x_9/n674 ) );
  NR2D0 U2222 ( .A1(n1802), .A2(n1822), .ZN(n1804) );
  OAI22D0 U2223 ( .A1(n1807), .A2(n1826), .B1(n1812), .B2(n1824), .ZN(n1803)
         );
  AOI211D0 U2224 ( .A1(n1805), .A2(n1830), .B(n1804), .C(n1803), .ZN(n1806) );
  MUX2ND0 U2225 ( .I0(R[5]), .I1(\mult_x_9/n660 ), .S(n1806), .ZN(
        \mult_x_9/n675 ) );
  NR2D0 U2226 ( .A1(n1807), .A2(n1822), .ZN(n1809) );
  OAI22D0 U2227 ( .A1(n1812), .A2(n1826), .B1(n1817), .B2(n1824), .ZN(n1808)
         );
  AOI211D0 U2228 ( .A1(n1810), .A2(n1830), .B(n1809), .C(n1808), .ZN(n1811) );
  MUX2ND0 U2229 ( .I0(R[5]), .I1(\mult_x_9/n660 ), .S(n1811), .ZN(
        \mult_x_9/n676 ) );
  NR2D0 U2230 ( .A1(n1812), .A2(n1822), .ZN(n1814) );
  OAI22D0 U2231 ( .A1(n1817), .A2(n1826), .B1(n1823), .B2(n1824), .ZN(n1813)
         );
  AOI211D0 U2232 ( .A1(n1815), .A2(n1830), .B(n1814), .C(n1813), .ZN(n1816) );
  MUX2ND0 U2233 ( .I0(R[5]), .I1(\mult_x_9/n660 ), .S(n1816), .ZN(
        \mult_x_9/n677 ) );
  NR2D0 U2234 ( .A1(n1817), .A2(n1822), .ZN(n1819) );
  OAI22D0 U2235 ( .A1(n1823), .A2(n1826), .B1(n1827), .B2(n1824), .ZN(n1818)
         );
  AOI211D0 U2236 ( .A1(n1820), .A2(n1830), .B(n1819), .C(n1818), .ZN(n1821) );
  MUX2ND0 U2237 ( .I0(R[5]), .I1(\mult_x_9/n660 ), .S(n1821), .ZN(
        \mult_x_9/n678 ) );
  NR2D0 U2238 ( .A1(n1823), .A2(n1822), .ZN(n1829) );
  OAI22D0 U2239 ( .A1(n1827), .A2(n1826), .B1(n1825), .B2(n1824), .ZN(n1828)
         );
  AOI211D0 U2240 ( .A1(n1831), .A2(n1830), .B(n1829), .C(n1828), .ZN(n1832) );
  MUX2ND0 U2241 ( .I0(R[5]), .I1(\mult_x_9/n660 ), .S(n1832), .ZN(
        \mult_x_9/n679 ) );
  FA1D0 U2242 ( .A(n2028), .B(\mult_x_13/n203 ), .CI(n1833), .CO(
        \mult_x_13/n188 ), .S(\mult_x_13/n197 ) );
  CKND2D0 U2243 ( .A1(R_lat_mag[17]), .A2(\mult_x_13/n382 ), .ZN(n1834) );
  MUX2ND0 U2244 ( .I0(n1836), .I1(n1835), .S(n1834), .ZN(\mult_x_13/n374 ) );
  CKND2D0 U2245 ( .A1(R_lat_mag[11]), .A2(\mult_x_13/n418 ), .ZN(n1837) );
  MUX2ND0 U2246 ( .I0(n1839), .I1(n1838), .S(n1837), .ZN(\mult_x_13/n413 ) );
  OAI222D0 U2247 ( .A1(n1844), .A2(n1843), .B1(n1842), .B2(n1841), .C1(n2174), 
        .C2(n1840), .ZN(\mult_x_13/n528 ) );
  NR2D0 U2248 ( .A1(n2185), .A2(n1893), .ZN(n1846) );
  OAI22D0 U2249 ( .A1(n2187), .A2(n1895), .B1(n2099), .B2(n1894), .ZN(n1845)
         );
  AOI211D0 U2250 ( .A1(n1898), .A2(n2190), .B(n1846), .C(n1845), .ZN(n1847) );
  MUX2ND0 U2251 ( .I0(R_lat_mag[20]), .I1(n1900), .S(n1847), .ZN(
        \mult_x_13/n533 ) );
  NR2D0 U2252 ( .A1(n2187), .A2(n1893), .ZN(n1849) );
  OAI22D0 U2253 ( .A1(n2099), .A2(n1895), .B1(n2103), .B2(n1894), .ZN(n1848)
         );
  AOI211D0 U2254 ( .A1(n1898), .A2(n2194), .B(n1849), .C(n1848), .ZN(n1850) );
  MUX2ND0 U2255 ( .I0(R_lat_mag[20]), .I1(n1900), .S(n1850), .ZN(
        \mult_x_13/n534 ) );
  NR2D0 U2256 ( .A1(n2099), .A2(n1893), .ZN(n1852) );
  OAI22D0 U2257 ( .A1(n2103), .A2(n1895), .B1(n2107), .B2(n1894), .ZN(n1851)
         );
  AOI211D0 U2258 ( .A1(n1898), .A2(n2198), .B(n1852), .C(n1851), .ZN(n1853) );
  MUX2ND0 U2259 ( .I0(R_lat_mag[20]), .I1(n1900), .S(n1853), .ZN(
        \mult_x_13/n535 ) );
  NR2D0 U2260 ( .A1(n2103), .A2(n1893), .ZN(n1855) );
  OAI22D0 U2261 ( .A1(n2107), .A2(n1895), .B1(n2111), .B2(n1894), .ZN(n1854)
         );
  AOI211D0 U2262 ( .A1(n1898), .A2(n2202), .B(n1855), .C(n1854), .ZN(n1856) );
  MUX2ND0 U2263 ( .I0(R_lat_mag[20]), .I1(n1900), .S(n1856), .ZN(
        \mult_x_13/n536 ) );
  NR2D0 U2264 ( .A1(n2107), .A2(n1893), .ZN(n1858) );
  OAI22D0 U2265 ( .A1(n2111), .A2(n1895), .B1(n2115), .B2(n1894), .ZN(n1857)
         );
  AOI211D0 U2266 ( .A1(n1898), .A2(n2206), .B(n1858), .C(n1857), .ZN(n1859) );
  MUX2ND0 U2267 ( .I0(R_lat_mag[20]), .I1(n1900), .S(n1859), .ZN(
        \mult_x_13/n537 ) );
  NR2D0 U2268 ( .A1(n2115), .A2(n1893), .ZN(n1861) );
  OAI22D0 U2269 ( .A1(n2119), .A2(n1895), .B1(n2123), .B2(n1894), .ZN(n1860)
         );
  AOI211D0 U2270 ( .A1(n1898), .A2(n2214), .B(n1861), .C(n1860), .ZN(n1862) );
  MUX2ND0 U2271 ( .I0(R_lat_mag[20]), .I1(n1900), .S(n1862), .ZN(
        \mult_x_13/n539 ) );
  OAI22D0 U2272 ( .A1(n2119), .A2(n1893), .B1(n2127), .B2(n1894), .ZN(n1863)
         );
  AOI211D0 U2273 ( .A1(n1898), .A2(n2218), .B(n1864), .C(n1863), .ZN(n1865) );
  MUX2ND0 U2274 ( .I0(R_lat_mag[20]), .I1(n1900), .S(n1865), .ZN(
        \mult_x_13/n540 ) );
  NR2D0 U2275 ( .A1(n2127), .A2(n1895), .ZN(n1867) );
  OAI22D0 U2276 ( .A1(n2123), .A2(n1893), .B1(n2131), .B2(n1894), .ZN(n1866)
         );
  AOI211D0 U2277 ( .A1(n1898), .A2(n2222), .B(n1867), .C(n1866), .ZN(n1868) );
  MUX2ND0 U2278 ( .I0(R_lat_mag[20]), .I1(n1900), .S(n1868), .ZN(
        \mult_x_13/n541 ) );
  NR2D0 U2279 ( .A1(n2127), .A2(n1893), .ZN(n1870) );
  OAI22D0 U2280 ( .A1(n2131), .A2(n1895), .B1(n2135), .B2(n1894), .ZN(n1869)
         );
  AOI211D0 U2281 ( .A1(n1898), .A2(n2226), .B(n1870), .C(n1869), .ZN(n1871) );
  MUX2ND0 U2282 ( .I0(R_lat_mag[20]), .I1(n1900), .S(n1871), .ZN(
        \mult_x_13/n542 ) );
  NR2D0 U2283 ( .A1(n2139), .A2(n1893), .ZN(n1873) );
  OAI22D0 U2284 ( .A1(n2147), .A2(n1894), .B1(n2143), .B2(n1895), .ZN(n1872)
         );
  AOI211D0 U2285 ( .A1(n1898), .A2(n2238), .B(n1873), .C(n1872), .ZN(n1874) );
  MUX2ND0 U2286 ( .I0(R_lat_mag[20]), .I1(n1900), .S(n1874), .ZN(
        \mult_x_13/n545 ) );
  NR2D0 U2287 ( .A1(n2143), .A2(n1893), .ZN(n1876) );
  OAI22D0 U2288 ( .A1(n2151), .A2(n1894), .B1(n2147), .B2(n1895), .ZN(n1875)
         );
  AOI211D0 U2289 ( .A1(n1898), .A2(n2242), .B(n1876), .C(n1875), .ZN(n1877) );
  MUX2ND0 U2290 ( .I0(R_lat_mag[20]), .I1(n1900), .S(n1877), .ZN(
        \mult_x_13/n546 ) );
  NR2D0 U2291 ( .A1(n2147), .A2(n1893), .ZN(n1879) );
  OAI22D0 U2292 ( .A1(n2155), .A2(n1894), .B1(n2151), .B2(n1895), .ZN(n1878)
         );
  AOI211D0 U2293 ( .A1(n1898), .A2(n2246), .B(n1879), .C(n1878), .ZN(n1880) );
  MUX2ND0 U2294 ( .I0(R_lat_mag[20]), .I1(n1900), .S(n1880), .ZN(
        \mult_x_13/n547 ) );
  NR2D0 U2295 ( .A1(n2151), .A2(n1893), .ZN(n1882) );
  OAI22D0 U2296 ( .A1(n2159), .A2(n1894), .B1(n2155), .B2(n1895), .ZN(n1881)
         );
  AOI211D0 U2297 ( .A1(n1898), .A2(n2250), .B(n1882), .C(n1881), .ZN(n1883) );
  MUX2ND0 U2298 ( .I0(R_lat_mag[20]), .I1(n1900), .S(n1883), .ZN(
        \mult_x_13/n548 ) );
  NR2D0 U2299 ( .A1(n2155), .A2(n1893), .ZN(n1885) );
  OAI22D0 U2300 ( .A1(n2164), .A2(n1894), .B1(n2159), .B2(n1895), .ZN(n1884)
         );
  AOI211D0 U2301 ( .A1(n1898), .A2(n2254), .B(n1885), .C(n1884), .ZN(n1886) );
  MUX2ND0 U2302 ( .I0(R_lat_mag[20]), .I1(n1900), .S(n1886), .ZN(
        \mult_x_13/n549 ) );
  NR2D0 U2303 ( .A1(n2159), .A2(n1893), .ZN(n1888) );
  OAI22D0 U2304 ( .A1(n2172), .A2(n1894), .B1(n2164), .B2(n1895), .ZN(n1887)
         );
  AOI211D0 U2305 ( .A1(n1898), .A2(n2162), .B(n1888), .C(n1887), .ZN(n1889) );
  MUX2ND0 U2306 ( .I0(R_lat_mag[20]), .I1(n1900), .S(n1889), .ZN(
        \mult_x_13/n550 ) );
  NR2D0 U2307 ( .A1(n2164), .A2(n1893), .ZN(n1891) );
  OAI22D0 U2308 ( .A1(n2170), .A2(n1894), .B1(n2172), .B2(n1895), .ZN(n1890)
         );
  AOI211D0 U2309 ( .A1(n1898), .A2(n2167), .B(n1891), .C(n1890), .ZN(n1892) );
  MUX2ND0 U2310 ( .I0(R_lat_mag[20]), .I1(n1900), .S(n1892), .ZN(
        \mult_x_13/n551 ) );
  OAI22D0 U2311 ( .A1(n2170), .A2(n1895), .B1(n2174), .B2(n1894), .ZN(n1896)
         );
  AOI211D0 U2312 ( .A1(n1898), .A2(n2177), .B(n1897), .C(n1896), .ZN(n1899) );
  MUX2ND0 U2313 ( .I0(R_lat_mag[20]), .I1(n1900), .S(n1899), .ZN(
        \mult_x_13/n552 ) );
  AOI22D0 U2314 ( .A1(inv_Q_mag[22]), .A2(n1955), .B1(n2181), .B2(n1954), .ZN(
        n1901) );
  MUX2ND0 U2315 ( .I0(R_lat_mag[17]), .I1(\mult_x_13/n556 ), .S(n1901), .ZN(
        \mult_x_13/n557 ) );
  INVD0 U2316 ( .I(n1957), .ZN(n1903) );
  OAI222D0 U2317 ( .A1(n1904), .A2(n2187), .B1(n1903), .B2(n2185), .C1(n2184), 
        .C2(n1902), .ZN(n1905) );
  MUX2ND0 U2318 ( .I0(\mult_x_13/n556 ), .I1(R_lat_mag[17]), .S(n1905), .ZN(
        \mult_x_13/n558 ) );
  AOI22D0 U2319 ( .A1(inv_Q_mag[20]), .A2(n1955), .B1(n2190), .B2(n1954), .ZN(
        n1907) );
  AOI22D0 U2320 ( .A1(inv_Q_mag[22]), .A2(n1956), .B1(inv_Q_mag[21]), .B2(
        n1957), .ZN(n1906) );
  CKND2D0 U2321 ( .A1(n1907), .A2(n1906), .ZN(n1908) );
  MUX2ND0 U2322 ( .I0(\mult_x_13/n556 ), .I1(R_lat_mag[17]), .S(n1908), .ZN(
        \mult_x_13/n559 ) );
  AOI22D0 U2323 ( .A1(inv_Q_mag[19]), .A2(n1955), .B1(n2194), .B2(n1954), .ZN(
        n1910) );
  AOI22D0 U2324 ( .A1(inv_Q_mag[21]), .A2(n1956), .B1(inv_Q_mag[20]), .B2(
        n1957), .ZN(n1909) );
  CKND2D0 U2325 ( .A1(n1910), .A2(n1909), .ZN(n1911) );
  MUX2ND0 U2326 ( .I0(\mult_x_13/n556 ), .I1(R_lat_mag[17]), .S(n1911), .ZN(
        \mult_x_13/n560 ) );
  AOI22D0 U2327 ( .A1(inv_Q_mag[18]), .A2(n1955), .B1(n2198), .B2(n1954), .ZN(
        n1913) );
  AOI22D0 U2328 ( .A1(inv_Q_mag[20]), .A2(n1956), .B1(inv_Q_mag[19]), .B2(
        n1957), .ZN(n1912) );
  MUX2ND0 U2329 ( .I0(\mult_x_13/n556 ), .I1(R_lat_mag[17]), .S(n1914), .ZN(
        \mult_x_13/n561 ) );
  AOI22D0 U2330 ( .A1(inv_Q_mag[17]), .A2(n1955), .B1(n2202), .B2(n1954), .ZN(
        n1916) );
  AOI22D0 U2331 ( .A1(inv_Q_mag[19]), .A2(n1956), .B1(inv_Q_mag[18]), .B2(
        n1957), .ZN(n1915) );
  CKND2D0 U2332 ( .A1(n1916), .A2(n1915), .ZN(n1917) );
  MUX2ND0 U2333 ( .I0(\mult_x_13/n556 ), .I1(R_lat_mag[17]), .S(n1917), .ZN(
        \mult_x_13/n562 ) );
  AOI22D0 U2334 ( .A1(inv_Q_mag[16]), .A2(n1955), .B1(n2206), .B2(n1954), .ZN(
        n1919) );
  AOI22D0 U2335 ( .A1(inv_Q_mag[18]), .A2(n1956), .B1(inv_Q_mag[17]), .B2(
        n1957), .ZN(n1918) );
  CKND2D0 U2336 ( .A1(n1919), .A2(n1918), .ZN(n1920) );
  MUX2ND0 U2337 ( .I0(\mult_x_13/n556 ), .I1(R_lat_mag[17]), .S(n1920), .ZN(
        \mult_x_13/n563 ) );
  AOI22D0 U2338 ( .A1(inv_Q_mag[17]), .A2(n1956), .B1(inv_Q_mag[16]), .B2(
        n1957), .ZN(n1921) );
  CKND2D0 U2339 ( .A1(n1922), .A2(n1921), .ZN(n1923) );
  MUX2ND0 U2340 ( .I0(\mult_x_13/n556 ), .I1(R_lat_mag[17]), .S(n1923), .ZN(
        \mult_x_13/n564 ) );
  AOI22D0 U2341 ( .A1(inv_Q_mag[14]), .A2(n1955), .B1(n2214), .B2(n1954), .ZN(
        n1925) );
  AOI22D0 U2342 ( .A1(inv_Q_mag[16]), .A2(n1956), .B1(inv_Q_mag[15]), .B2(
        n1957), .ZN(n1924) );
  CKND2D0 U2343 ( .A1(n1925), .A2(n1924), .ZN(n1926) );
  MUX2ND0 U2344 ( .I0(\mult_x_13/n556 ), .I1(R_lat_mag[17]), .S(n1926), .ZN(
        \mult_x_13/n565 ) );
  AOI22D0 U2345 ( .A1(inv_Q_mag[15]), .A2(n1956), .B1(n2218), .B2(n1954), .ZN(
        n1928) );
  CKND2D0 U2346 ( .A1(n1928), .A2(n1927), .ZN(n1929) );
  MUX2ND0 U2347 ( .I0(\mult_x_13/n556 ), .I1(R_lat_mag[17]), .S(n1929), .ZN(
        \mult_x_13/n566 ) );
  AOI22D0 U2348 ( .A1(inv_Q_mag[14]), .A2(n1956), .B1(n2222), .B2(n1954), .ZN(
        n1931) );
  AOI22D0 U2349 ( .A1(inv_Q_mag[13]), .A2(n1957), .B1(inv_Q_mag[12]), .B2(
        n1955), .ZN(n1930) );
  MUX2ND0 U2350 ( .I0(\mult_x_13/n556 ), .I1(R_lat_mag[17]), .S(n1932), .ZN(
        \mult_x_13/n567 ) );
  AOI22D0 U2351 ( .A1(inv_Q_mag[11]), .A2(n1955), .B1(n2226), .B2(n1954), .ZN(
        n1934) );
  AOI22D0 U2352 ( .A1(inv_Q_mag[13]), .A2(n1956), .B1(inv_Q_mag[12]), .B2(
        n1957), .ZN(n1933) );
  CKND2D0 U2353 ( .A1(n1934), .A2(n1933), .ZN(n1935) );
  MUX2ND0 U2354 ( .I0(\mult_x_13/n556 ), .I1(R_lat_mag[17]), .S(n1935), .ZN(
        \mult_x_13/n568 ) );
  AOI22D0 U2355 ( .A1(inv_Q_mag[10]), .A2(n1955), .B1(n2230), .B2(n1954), .ZN(
        n1937) );
  AOI22D0 U2356 ( .A1(inv_Q_mag[12]), .A2(n1956), .B1(inv_Q_mag[11]), .B2(
        n1957), .ZN(n1936) );
  CKND2D0 U2357 ( .A1(n1937), .A2(n1936), .ZN(n1938) );
  MUX2ND0 U2358 ( .I0(\mult_x_13/n556 ), .I1(R_lat_mag[17]), .S(n1938), .ZN(
        \mult_x_13/n569 ) );
  AOI22D0 U2359 ( .A1(inv_Q_mag[9]), .A2(n1955), .B1(n2234), .B2(n1954), .ZN(
        n1940) );
  AOI22D0 U2360 ( .A1(inv_Q_mag[10]), .A2(n1957), .B1(inv_Q_mag[11]), .B2(
        n1956), .ZN(n1939) );
  CKND2D0 U2361 ( .A1(n1940), .A2(n1939), .ZN(n1941) );
  MUX2ND0 U2362 ( .I0(\mult_x_13/n556 ), .I1(R_lat_mag[17]), .S(n1941), .ZN(
        \mult_x_13/n570 ) );
  AOI22D0 U2363 ( .A1(inv_Q_mag[8]), .A2(n1955), .B1(n2238), .B2(n1954), .ZN(
        n1943) );
  AOI22D0 U2364 ( .A1(inv_Q_mag[9]), .A2(n1957), .B1(inv_Q_mag[10]), .B2(n1956), .ZN(n1942) );
  CKND2D0 U2365 ( .A1(n1943), .A2(n1942), .ZN(n1944) );
  MUX2ND0 U2366 ( .I0(\mult_x_13/n556 ), .I1(R_lat_mag[17]), .S(n1944), .ZN(
        \mult_x_13/n571 ) );
  AOI22D0 U2367 ( .A1(inv_Q_mag[8]), .A2(n1957), .B1(inv_Q_mag[9]), .B2(n1956), 
        .ZN(n1945) );
  CKND2D0 U2368 ( .A1(n1946), .A2(n1945), .ZN(n1947) );
  MUX2ND0 U2369 ( .I0(\mult_x_13/n556 ), .I1(R_lat_mag[17]), .S(n1947), .ZN(
        \mult_x_13/n572 ) );
  AOI22D0 U2370 ( .A1(inv_Q_mag[6]), .A2(n1955), .B1(n2246), .B2(n1954), .ZN(
        n1949) );
  AOI22D0 U2371 ( .A1(inv_Q_mag[7]), .A2(n1957), .B1(inv_Q_mag[8]), .B2(n1956), 
        .ZN(n1948) );
  CKND2D0 U2372 ( .A1(n1949), .A2(n1948), .ZN(n1950) );
  MUX2ND0 U2373 ( .I0(\mult_x_13/n556 ), .I1(R_lat_mag[17]), .S(n1950), .ZN(
        \mult_x_13/n573 ) );
  AOI22D0 U2374 ( .A1(inv_Q_mag[5]), .A2(n1955), .B1(n2250), .B2(n1954), .ZN(
        n1952) );
  AOI22D0 U2375 ( .A1(inv_Q_mag[6]), .A2(n1957), .B1(inv_Q_mag[7]), .B2(n1956), 
        .ZN(n1951) );
  MUX2ND0 U2376 ( .I0(\mult_x_13/n556 ), .I1(R_lat_mag[17]), .S(n1953), .ZN(
        \mult_x_13/n574 ) );
  AOI22D0 U2377 ( .A1(inv_Q_mag[4]), .A2(n1955), .B1(n2254), .B2(n1954), .ZN(
        n1959) );
  AOI22D0 U2378 ( .A1(inv_Q_mag[5]), .A2(n1957), .B1(inv_Q_mag[6]), .B2(n1956), 
        .ZN(n1958) );
  CKND2D0 U2379 ( .A1(n1959), .A2(n1958), .ZN(n1960) );
  MUX2ND0 U2380 ( .I0(\mult_x_13/n556 ), .I1(R_lat_mag[17]), .S(n1960), .ZN(
        \mult_x_13/n575 ) );
  OAI22D0 U2381 ( .A1(n2185), .A2(n2023), .B1(n2089), .B2(n1962), .ZN(n1961)
         );
  MUX2ND0 U2382 ( .I0(n2028), .I1(R_lat_mag[14]), .S(n1961), .ZN(
        \mult_x_13/n583 ) );
  OAI222D0 U2383 ( .A1(n2023), .A2(n2187), .B1(n2021), .B2(n2185), .C1(n2184), 
        .C2(n1962), .ZN(n1963) );
  MUX2ND0 U2384 ( .I0(n2028), .I1(R_lat_mag[14]), .S(n1963), .ZN(
        \mult_x_13/n584 ) );
  NR2D0 U2385 ( .A1(n2187), .A2(n2021), .ZN(n1965) );
  AOI211D0 U2386 ( .A1(n2026), .A2(n2190), .B(n1965), .C(n1964), .ZN(n1966) );
  MUX2ND0 U2387 ( .I0(R_lat_mag[14]), .I1(n2028), .S(n1966), .ZN(
        \mult_x_13/n585 ) );
  NR2D0 U2388 ( .A1(n2099), .A2(n2021), .ZN(n1968) );
  OAI22D0 U2389 ( .A1(n2187), .A2(n2022), .B1(n2103), .B2(n2023), .ZN(n1967)
         );
  AOI211D0 U2390 ( .A1(n2026), .A2(n2194), .B(n1968), .C(n1967), .ZN(n1969) );
  MUX2ND0 U2391 ( .I0(R_lat_mag[14]), .I1(n2028), .S(n1969), .ZN(
        \mult_x_13/n586 ) );
  NR2D0 U2392 ( .A1(n2103), .A2(n2021), .ZN(n1971) );
  OAI22D0 U2393 ( .A1(n2099), .A2(n2022), .B1(n2107), .B2(n2023), .ZN(n1970)
         );
  MUX2ND0 U2394 ( .I0(R_lat_mag[14]), .I1(n2028), .S(n1972), .ZN(
        \mult_x_13/n587 ) );
  NR2D0 U2395 ( .A1(n2107), .A2(n2021), .ZN(n1974) );
  AOI211D0 U2396 ( .A1(n2026), .A2(n2202), .B(n1974), .C(n1973), .ZN(n1975) );
  MUX2ND0 U2397 ( .I0(R_lat_mag[14]), .I1(n2028), .S(n1975), .ZN(
        \mult_x_13/n588 ) );
  NR2D0 U2398 ( .A1(n2111), .A2(n2021), .ZN(n1977) );
  OAI22D0 U2399 ( .A1(n2107), .A2(n2022), .B1(n2115), .B2(n2023), .ZN(n1976)
         );
  AOI211D0 U2400 ( .A1(n2026), .A2(n2206), .B(n1977), .C(n1976), .ZN(n1978) );
  MUX2ND0 U2401 ( .I0(R_lat_mag[14]), .I1(n2028), .S(n1978), .ZN(
        \mult_x_13/n589 ) );
  NR2D0 U2402 ( .A1(n2115), .A2(n2021), .ZN(n1980) );
  OAI22D0 U2403 ( .A1(n2111), .A2(n2022), .B1(n2119), .B2(n2023), .ZN(n1979)
         );
  AOI211D0 U2404 ( .A1(n2026), .A2(n2210), .B(n1980), .C(n1979), .ZN(n1981) );
  MUX2ND0 U2405 ( .I0(R_lat_mag[14]), .I1(n2028), .S(n1981), .ZN(
        \mult_x_13/n590 ) );
  NR2D0 U2406 ( .A1(n2119), .A2(n2021), .ZN(n1983) );
  OAI22D0 U2407 ( .A1(n2115), .A2(n2022), .B1(n2123), .B2(n2023), .ZN(n1982)
         );
  AOI211D0 U2408 ( .A1(n2026), .A2(n2214), .B(n1983), .C(n1982), .ZN(n1984) );
  MUX2ND0 U2409 ( .I0(R_lat_mag[14]), .I1(n2028), .S(n1984), .ZN(
        \mult_x_13/n591 ) );
  NR2D0 U2410 ( .A1(n2127), .A2(n2023), .ZN(n1986) );
  AOI211D0 U2411 ( .A1(n2026), .A2(n2218), .B(n1986), .C(n1985), .ZN(n1987) );
  MUX2ND0 U2412 ( .I0(R_lat_mag[14]), .I1(n2028), .S(n1987), .ZN(
        \mult_x_13/n592 ) );
  NR2D0 U2413 ( .A1(n2131), .A2(n2023), .ZN(n1989) );
  OAI22D0 U2414 ( .A1(n2123), .A2(n2022), .B1(n2127), .B2(n2021), .ZN(n1988)
         );
  AOI211D0 U2415 ( .A1(n2026), .A2(n2222), .B(n1989), .C(n1988), .ZN(n1990) );
  MUX2ND0 U2416 ( .I0(R_lat_mag[14]), .I1(n2028), .S(n1990), .ZN(
        \mult_x_13/n593 ) );
  NR2D0 U2417 ( .A1(n2131), .A2(n2021), .ZN(n1992) );
  OAI22D0 U2418 ( .A1(n2127), .A2(n2022), .B1(n2135), .B2(n2023), .ZN(n1991)
         );
  AOI211D0 U2419 ( .A1(n2026), .A2(n2226), .B(n1992), .C(n1991), .ZN(n1993) );
  MUX2ND0 U2420 ( .I0(R_lat_mag[14]), .I1(n2028), .S(n1993), .ZN(
        \mult_x_13/n594 ) );
  NR2D0 U2421 ( .A1(n2135), .A2(n2021), .ZN(n1995) );
  OAI22D0 U2422 ( .A1(n2131), .A2(n2022), .B1(n2139), .B2(n2023), .ZN(n1994)
         );
  AOI211D0 U2423 ( .A1(n2026), .A2(n2230), .B(n1995), .C(n1994), .ZN(n1996) );
  MUX2ND0 U2424 ( .I0(R_lat_mag[14]), .I1(n2028), .S(n1996), .ZN(
        \mult_x_13/n595 ) );
  NR2D0 U2425 ( .A1(n2139), .A2(n2021), .ZN(n1998) );
  OAI22D0 U2426 ( .A1(n2143), .A2(n2023), .B1(n2135), .B2(n2022), .ZN(n1997)
         );
  AOI211D0 U2427 ( .A1(n2026), .A2(n2234), .B(n1998), .C(n1997), .ZN(n1999) );
  MUX2ND0 U2428 ( .I0(R_lat_mag[14]), .I1(n2028), .S(n1999), .ZN(
        \mult_x_13/n596 ) );
  NR2D0 U2429 ( .A1(n2143), .A2(n2021), .ZN(n2001) );
  OAI22D0 U2430 ( .A1(n2147), .A2(n2023), .B1(n2139), .B2(n2022), .ZN(n2000)
         );
  AOI211D0 U2431 ( .A1(n2026), .A2(n2238), .B(n2001), .C(n2000), .ZN(n2002) );
  MUX2ND0 U2432 ( .I0(R_lat_mag[14]), .I1(n2028), .S(n2002), .ZN(
        \mult_x_13/n597 ) );
  NR2D0 U2433 ( .A1(n2147), .A2(n2021), .ZN(n2004) );
  OAI22D0 U2434 ( .A1(n2151), .A2(n2023), .B1(n2143), .B2(n2022), .ZN(n2003)
         );
  AOI211D0 U2435 ( .A1(n2026), .A2(n2242), .B(n2004), .C(n2003), .ZN(n2005) );
  MUX2ND0 U2436 ( .I0(R_lat_mag[14]), .I1(n2028), .S(n2005), .ZN(
        \mult_x_13/n598 ) );
  NR2D0 U2437 ( .A1(n2151), .A2(n2021), .ZN(n2007) );
  OAI22D0 U2438 ( .A1(n2155), .A2(n2023), .B1(n2147), .B2(n2022), .ZN(n2006)
         );
  AOI211D0 U2439 ( .A1(n2026), .A2(n2246), .B(n2007), .C(n2006), .ZN(n2008) );
  MUX2ND0 U2440 ( .I0(R_lat_mag[14]), .I1(n2028), .S(n2008), .ZN(
        \mult_x_13/n599 ) );
  NR2D0 U2441 ( .A1(n2155), .A2(n2021), .ZN(n2010) );
  OAI22D0 U2442 ( .A1(n2159), .A2(n2023), .B1(n2151), .B2(n2022), .ZN(n2009)
         );
  AOI211D0 U2443 ( .A1(n2026), .A2(n2250), .B(n2010), .C(n2009), .ZN(n2011) );
  MUX2ND0 U2444 ( .I0(R_lat_mag[14]), .I1(n2028), .S(n2011), .ZN(
        \mult_x_13/n600 ) );
  NR2D0 U2445 ( .A1(n2159), .A2(n2021), .ZN(n2013) );
  AOI211D0 U2446 ( .A1(n2026), .A2(n2254), .B(n2013), .C(n2012), .ZN(n2014) );
  MUX2ND0 U2447 ( .I0(R_lat_mag[14]), .I1(n2028), .S(n2014), .ZN(
        \mult_x_13/n601 ) );
  NR2D0 U2448 ( .A1(n2164), .A2(n2021), .ZN(n2016) );
  OAI22D0 U2449 ( .A1(n2172), .A2(n2023), .B1(n2159), .B2(n2022), .ZN(n2015)
         );
  AOI211D0 U2450 ( .A1(n2026), .A2(n2162), .B(n2016), .C(n2015), .ZN(n2017) );
  MUX2ND0 U2451 ( .I0(R_lat_mag[14]), .I1(n2028), .S(n2017), .ZN(
        \mult_x_13/n602 ) );
  NR2D0 U2452 ( .A1(n2172), .A2(n2021), .ZN(n2019) );
  OAI22D0 U2453 ( .A1(n2170), .A2(n2023), .B1(n2164), .B2(n2022), .ZN(n2018)
         );
  AOI211D0 U2454 ( .A1(n2026), .A2(n2167), .B(n2019), .C(n2018), .ZN(n2020) );
  MUX2ND0 U2455 ( .I0(R_lat_mag[14]), .I1(n2028), .S(n2020), .ZN(
        \mult_x_13/n603 ) );
  NR2D0 U2456 ( .A1(n2170), .A2(n2021), .ZN(n2025) );
  OAI22D0 U2457 ( .A1(n2174), .A2(n2023), .B1(n2172), .B2(n2022), .ZN(n2024)
         );
  AOI211D0 U2458 ( .A1(n2026), .A2(n2177), .B(n2025), .C(n2024), .ZN(n2027) );
  MUX2ND0 U2459 ( .I0(R_lat_mag[14]), .I1(n2028), .S(n2027), .ZN(
        \mult_x_13/n604 ) );
  AOI22D0 U2460 ( .A1(inv_Q_mag[22]), .A2(n2083), .B1(n2181), .B2(n2082), .ZN(
        n2029) );
  MUX2ND0 U2461 ( .I0(R_lat_mag[11]), .I1(\mult_x_13/n608 ), .S(n2029), .ZN(
        \mult_x_13/n609 ) );
  INVD0 U2462 ( .I(n2085), .ZN(n2031) );
  OAI222D0 U2463 ( .A1(n2032), .A2(n2187), .B1(n2031), .B2(n2185), .C1(n2184), 
        .C2(n2030), .ZN(n2033) );
  MUX2ND0 U2464 ( .I0(\mult_x_13/n608 ), .I1(R_lat_mag[11]), .S(n2033), .ZN(
        \mult_x_13/n610 ) );
  AOI22D0 U2465 ( .A1(inv_Q_mag[20]), .A2(n2083), .B1(n2190), .B2(n2082), .ZN(
        n2035) );
  AOI22D0 U2466 ( .A1(inv_Q_mag[22]), .A2(n2084), .B1(inv_Q_mag[21]), .B2(
        n2085), .ZN(n2034) );
  MUX2ND0 U2467 ( .I0(\mult_x_13/n608 ), .I1(R_lat_mag[11]), .S(n2036), .ZN(
        \mult_x_13/n611 ) );
  AOI22D0 U2468 ( .A1(inv_Q_mag[19]), .A2(n2083), .B1(n2194), .B2(n2082), .ZN(
        n2038) );
  AOI22D0 U2469 ( .A1(inv_Q_mag[21]), .A2(n2084), .B1(inv_Q_mag[20]), .B2(
        n2085), .ZN(n2037) );
  CKND2D0 U2470 ( .A1(n2038), .A2(n2037), .ZN(n2039) );
  MUX2ND0 U2471 ( .I0(\mult_x_13/n608 ), .I1(R_lat_mag[11]), .S(n2039), .ZN(
        \mult_x_13/n612 ) );
  AOI22D0 U2472 ( .A1(inv_Q_mag[18]), .A2(n2083), .B1(n2198), .B2(n2082), .ZN(
        n2041) );
  AOI22D0 U2473 ( .A1(inv_Q_mag[20]), .A2(n2084), .B1(inv_Q_mag[19]), .B2(
        n2085), .ZN(n2040) );
  MUX2ND0 U2474 ( .I0(\mult_x_13/n608 ), .I1(R_lat_mag[11]), .S(n2042), .ZN(
        \mult_x_13/n613 ) );
  AOI22D0 U2475 ( .A1(inv_Q_mag[17]), .A2(n2083), .B1(n2202), .B2(n2082), .ZN(
        n2044) );
  AOI22D0 U2476 ( .A1(inv_Q_mag[19]), .A2(n2084), .B1(inv_Q_mag[18]), .B2(
        n2085), .ZN(n2043) );
  CKND2D0 U2477 ( .A1(n2044), .A2(n2043), .ZN(n2045) );
  MUX2ND0 U2478 ( .I0(\mult_x_13/n608 ), .I1(R_lat_mag[11]), .S(n2045), .ZN(
        \mult_x_13/n614 ) );
  AOI22D0 U2479 ( .A1(inv_Q_mag[16]), .A2(n2083), .B1(n2206), .B2(n2082), .ZN(
        n2047) );
  AOI22D0 U2480 ( .A1(inv_Q_mag[18]), .A2(n2084), .B1(inv_Q_mag[17]), .B2(
        n2085), .ZN(n2046) );
  CKND2D0 U2481 ( .A1(n2047), .A2(n2046), .ZN(n2048) );
  MUX2ND0 U2482 ( .I0(\mult_x_13/n608 ), .I1(R_lat_mag[11]), .S(n2048), .ZN(
        \mult_x_13/n615 ) );
  AOI22D0 U2483 ( .A1(inv_Q_mag[15]), .A2(n2083), .B1(n2210), .B2(n2082), .ZN(
        n2050) );
  AOI22D0 U2484 ( .A1(inv_Q_mag[17]), .A2(n2084), .B1(inv_Q_mag[16]), .B2(
        n2085), .ZN(n2049) );
  CKND2D0 U2485 ( .A1(n2050), .A2(n2049), .ZN(n2051) );
  MUX2ND0 U2486 ( .I0(\mult_x_13/n608 ), .I1(R_lat_mag[11]), .S(n2051), .ZN(
        \mult_x_13/n616 ) );
  AOI22D0 U2487 ( .A1(inv_Q_mag[16]), .A2(n2084), .B1(inv_Q_mag[15]), .B2(
        n2085), .ZN(n2052) );
  CKND2D0 U2488 ( .A1(n2053), .A2(n2052), .ZN(n2054) );
  MUX2ND0 U2489 ( .I0(\mult_x_13/n608 ), .I1(R_lat_mag[11]), .S(n2054), .ZN(
        \mult_x_13/n617 ) );
  AOI22D0 U2490 ( .A1(inv_Q_mag[15]), .A2(n2084), .B1(n2218), .B2(n2082), .ZN(
        n2056) );
  AOI22D0 U2491 ( .A1(inv_Q_mag[14]), .A2(n2085), .B1(inv_Q_mag[13]), .B2(
        n2083), .ZN(n2055) );
  CKND2D0 U2492 ( .A1(n2056), .A2(n2055), .ZN(n2057) );
  MUX2ND0 U2493 ( .I0(\mult_x_13/n608 ), .I1(R_lat_mag[11]), .S(n2057), .ZN(
        \mult_x_13/n618 ) );
  AOI22D0 U2494 ( .A1(inv_Q_mag[14]), .A2(n2084), .B1(n2222), .B2(n2082), .ZN(
        n2059) );
  AOI22D0 U2495 ( .A1(inv_Q_mag[13]), .A2(n2085), .B1(inv_Q_mag[12]), .B2(
        n2083), .ZN(n2058) );
  CKND2D0 U2496 ( .A1(n2059), .A2(n2058), .ZN(n2060) );
  MUX2ND0 U2497 ( .I0(\mult_x_13/n608 ), .I1(R_lat_mag[11]), .S(n2060), .ZN(
        \mult_x_13/n619 ) );
  AOI22D0 U2498 ( .A1(inv_Q_mag[11]), .A2(n2083), .B1(n2226), .B2(n2082), .ZN(
        n2062) );
  AOI22D0 U2499 ( .A1(inv_Q_mag[13]), .A2(n2084), .B1(inv_Q_mag[12]), .B2(
        n2085), .ZN(n2061) );
  MUX2ND0 U2500 ( .I0(\mult_x_13/n608 ), .I1(R_lat_mag[11]), .S(n2063), .ZN(
        \mult_x_13/n620 ) );
  AOI22D0 U2501 ( .A1(inv_Q_mag[10]), .A2(n2083), .B1(n2230), .B2(n2082), .ZN(
        n2065) );
  AOI22D0 U2502 ( .A1(inv_Q_mag[12]), .A2(n2084), .B1(inv_Q_mag[11]), .B2(
        n2085), .ZN(n2064) );
  CKND2D0 U2503 ( .A1(n2065), .A2(n2064), .ZN(n2066) );
  MUX2ND0 U2504 ( .I0(\mult_x_13/n608 ), .I1(R_lat_mag[11]), .S(n2066), .ZN(
        \mult_x_13/n621 ) );
  AOI22D0 U2505 ( .A1(inv_Q_mag[10]), .A2(n2085), .B1(inv_Q_mag[11]), .B2(
        n2084), .ZN(n2067) );
  CKND2D0 U2506 ( .A1(n2068), .A2(n2067), .ZN(n2069) );
  MUX2ND0 U2507 ( .I0(\mult_x_13/n608 ), .I1(R_lat_mag[11]), .S(n2069), .ZN(
        \mult_x_13/n622 ) );
  AOI22D0 U2508 ( .A1(inv_Q_mag[8]), .A2(n2083), .B1(n2238), .B2(n2082), .ZN(
        n2071) );
  AOI22D0 U2509 ( .A1(inv_Q_mag[9]), .A2(n2085), .B1(inv_Q_mag[10]), .B2(n2084), .ZN(n2070) );
  CKND2D0 U2510 ( .A1(n2071), .A2(n2070), .ZN(n2072) );
  MUX2ND0 U2511 ( .I0(\mult_x_13/n608 ), .I1(R_lat_mag[11]), .S(n2072), .ZN(
        \mult_x_13/n623 ) );
  AOI22D0 U2512 ( .A1(inv_Q_mag[7]), .A2(n2083), .B1(n2242), .B2(n2082), .ZN(
        n2074) );
  AOI22D0 U2513 ( .A1(inv_Q_mag[8]), .A2(n2085), .B1(inv_Q_mag[9]), .B2(n2084), 
        .ZN(n2073) );
  CKND2D0 U2514 ( .A1(n2074), .A2(n2073), .ZN(n2075) );
  MUX2ND0 U2515 ( .I0(\mult_x_13/n608 ), .I1(R_lat_mag[11]), .S(n2075), .ZN(
        \mult_x_13/n624 ) );
  AOI22D0 U2516 ( .A1(inv_Q_mag[6]), .A2(n2083), .B1(n2246), .B2(n2082), .ZN(
        n2077) );
  AOI22D0 U2517 ( .A1(inv_Q_mag[7]), .A2(n2085), .B1(inv_Q_mag[8]), .B2(n2084), 
        .ZN(n2076) );
  MUX2ND0 U2518 ( .I0(\mult_x_13/n608 ), .I1(R_lat_mag[11]), .S(n2078), .ZN(
        \mult_x_13/n625 ) );
  AOI22D0 U2519 ( .A1(inv_Q_mag[6]), .A2(n2085), .B1(inv_Q_mag[7]), .B2(n2084), 
        .ZN(n2079) );
  CKND2D0 U2520 ( .A1(n2080), .A2(n2079), .ZN(n2081) );
  MUX2ND0 U2521 ( .I0(\mult_x_13/n608 ), .I1(R_lat_mag[11]), .S(n2081), .ZN(
        \mult_x_13/n626 ) );
  AOI22D0 U2522 ( .A1(inv_Q_mag[4]), .A2(n2083), .B1(n2254), .B2(n2082), .ZN(
        n2087) );
  AOI22D0 U2523 ( .A1(inv_Q_mag[5]), .A2(n2085), .B1(inv_Q_mag[6]), .B2(n2084), 
        .ZN(n2086) );
  CKND2D0 U2524 ( .A1(n2087), .A2(n2086), .ZN(n2088) );
  MUX2ND0 U2525 ( .I0(\mult_x_13/n608 ), .I1(R_lat_mag[11]), .S(n2088), .ZN(
        \mult_x_13/n627 ) );
  OAI22D0 U2526 ( .A1(n2185), .A2(n2173), .B1(n2089), .B2(n2091), .ZN(n2090)
         );
  MUX2ND0 U2527 ( .I0(n2180), .I1(R_lat_mag[8]), .S(n2090), .ZN(
        \mult_x_13/n635 ) );
  OAI222D0 U2528 ( .A1(n2173), .A2(n2187), .B1(n2169), .B2(n2185), .C1(n2184), 
        .C2(n2091), .ZN(n2092) );
  MUX2ND0 U2529 ( .I0(n2180), .I1(R_lat_mag[8]), .S(n2092), .ZN(
        \mult_x_13/n636 ) );
  NR2D0 U2530 ( .A1(n2187), .A2(n2169), .ZN(n2094) );
  OAI22D0 U2531 ( .A1(n2185), .A2(n2171), .B1(n2099), .B2(n2173), .ZN(n2093)
         );
  AOI211D0 U2532 ( .A1(n2178), .A2(n2190), .B(n2094), .C(n2093), .ZN(n2095) );
  MUX2ND0 U2533 ( .I0(R_lat_mag[8]), .I1(n2180), .S(n2095), .ZN(
        \mult_x_13/n637 ) );
  NR2D0 U2534 ( .A1(n2099), .A2(n2169), .ZN(n2097) );
  OAI22D0 U2535 ( .A1(n2187), .A2(n2171), .B1(n2103), .B2(n2173), .ZN(n2096)
         );
  AOI211D0 U2536 ( .A1(n2178), .A2(n2194), .B(n2097), .C(n2096), .ZN(n2098) );
  MUX2ND0 U2537 ( .I0(R_lat_mag[8]), .I1(n2180), .S(n2098), .ZN(
        \mult_x_13/n638 ) );
  NR2D0 U2538 ( .A1(n2103), .A2(n2169), .ZN(n2101) );
  OAI22D0 U2539 ( .A1(n2099), .A2(n2171), .B1(n2107), .B2(n2173), .ZN(n2100)
         );
  MUX2ND0 U2540 ( .I0(R_lat_mag[8]), .I1(n2180), .S(n2102), .ZN(
        \mult_x_13/n639 ) );
  NR2D0 U2541 ( .A1(n2107), .A2(n2169), .ZN(n2105) );
  OAI22D0 U2542 ( .A1(n2103), .A2(n2171), .B1(n2111), .B2(n2173), .ZN(n2104)
         );
  MUX2ND0 U2543 ( .I0(R_lat_mag[8]), .I1(n2180), .S(n2106), .ZN(
        \mult_x_13/n640 ) );
  NR2D0 U2544 ( .A1(n2111), .A2(n2169), .ZN(n2109) );
  OAI22D0 U2545 ( .A1(n2107), .A2(n2171), .B1(n2115), .B2(n2173), .ZN(n2108)
         );
  AOI211D0 U2546 ( .A1(n2178), .A2(n2206), .B(n2109), .C(n2108), .ZN(n2110) );
  MUX2ND0 U2547 ( .I0(R_lat_mag[8]), .I1(n2180), .S(n2110), .ZN(
        \mult_x_13/n641 ) );
  NR2D0 U2548 ( .A1(n2115), .A2(n2169), .ZN(n2113) );
  OAI22D0 U2549 ( .A1(n2111), .A2(n2171), .B1(n2119), .B2(n2173), .ZN(n2112)
         );
  AOI211D0 U2550 ( .A1(n2178), .A2(n2210), .B(n2113), .C(n2112), .ZN(n2114) );
  MUX2ND0 U2551 ( .I0(R_lat_mag[8]), .I1(n2180), .S(n2114), .ZN(
        \mult_x_13/n642 ) );
  NR2D0 U2552 ( .A1(n2119), .A2(n2169), .ZN(n2117) );
  OAI22D0 U2553 ( .A1(n2115), .A2(n2171), .B1(n2123), .B2(n2173), .ZN(n2116)
         );
  AOI211D0 U2554 ( .A1(n2178), .A2(n2214), .B(n2117), .C(n2116), .ZN(n2118) );
  MUX2ND0 U2555 ( .I0(R_lat_mag[8]), .I1(n2180), .S(n2118), .ZN(
        \mult_x_13/n643 ) );
  NR2D0 U2556 ( .A1(n2127), .A2(n2173), .ZN(n2121) );
  OAI22D0 U2557 ( .A1(n2119), .A2(n2171), .B1(n2123), .B2(n2169), .ZN(n2120)
         );
  AOI211D0 U2558 ( .A1(n2178), .A2(n2218), .B(n2121), .C(n2120), .ZN(n2122) );
  MUX2ND0 U2559 ( .I0(R_lat_mag[8]), .I1(n2180), .S(n2122), .ZN(
        \mult_x_13/n644 ) );
  NR2D0 U2560 ( .A1(n2131), .A2(n2173), .ZN(n2125) );
  OAI22D0 U2561 ( .A1(n2123), .A2(n2171), .B1(n2127), .B2(n2169), .ZN(n2124)
         );
  AOI211D0 U2562 ( .A1(n2178), .A2(n2222), .B(n2125), .C(n2124), .ZN(n2126) );
  MUX2ND0 U2563 ( .I0(R_lat_mag[8]), .I1(n2180), .S(n2126), .ZN(
        \mult_x_13/n645 ) );
  NR2D0 U2564 ( .A1(n2131), .A2(n2169), .ZN(n2129) );
  OAI22D0 U2565 ( .A1(n2127), .A2(n2171), .B1(n2135), .B2(n2173), .ZN(n2128)
         );
  AOI211D0 U2566 ( .A1(n2178), .A2(n2226), .B(n2129), .C(n2128), .ZN(n2130) );
  MUX2ND0 U2567 ( .I0(R_lat_mag[8]), .I1(n2180), .S(n2130), .ZN(
        \mult_x_13/n646 ) );
  NR2D0 U2568 ( .A1(n2135), .A2(n2169), .ZN(n2133) );
  OAI22D0 U2569 ( .A1(n2131), .A2(n2171), .B1(n2139), .B2(n2173), .ZN(n2132)
         );
  AOI211D0 U2570 ( .A1(n2178), .A2(n2230), .B(n2133), .C(n2132), .ZN(n2134) );
  MUX2ND0 U2571 ( .I0(R_lat_mag[8]), .I1(n2180), .S(n2134), .ZN(
        \mult_x_13/n647 ) );
  NR2D0 U2572 ( .A1(n2139), .A2(n2169), .ZN(n2137) );
  OAI22D0 U2573 ( .A1(n2143), .A2(n2173), .B1(n2135), .B2(n2171), .ZN(n2136)
         );
  AOI211D0 U2574 ( .A1(n2178), .A2(n2234), .B(n2137), .C(n2136), .ZN(n2138) );
  MUX2ND0 U2575 ( .I0(R_lat_mag[8]), .I1(n2180), .S(n2138), .ZN(
        \mult_x_13/n648 ) );
  NR2D0 U2576 ( .A1(n2143), .A2(n2169), .ZN(n2141) );
  OAI22D0 U2577 ( .A1(n2147), .A2(n2173), .B1(n2139), .B2(n2171), .ZN(n2140)
         );
  AOI211D0 U2578 ( .A1(n2178), .A2(n2238), .B(n2141), .C(n2140), .ZN(n2142) );
  MUX2ND0 U2579 ( .I0(R_lat_mag[8]), .I1(n2180), .S(n2142), .ZN(
        \mult_x_13/n649 ) );
  OAI22D0 U2580 ( .A1(n2151), .A2(n2173), .B1(n2143), .B2(n2171), .ZN(n2144)
         );
  AOI211D0 U2581 ( .A1(n2178), .A2(n2242), .B(n2145), .C(n2144), .ZN(n2146) );
  MUX2ND0 U2582 ( .I0(R_lat_mag[8]), .I1(n2180), .S(n2146), .ZN(
        \mult_x_13/n650 ) );
  NR2D0 U2583 ( .A1(n2151), .A2(n2169), .ZN(n2149) );
  OAI22D0 U2584 ( .A1(n2155), .A2(n2173), .B1(n2147), .B2(n2171), .ZN(n2148)
         );
  AOI211D0 U2585 ( .A1(n2178), .A2(n2246), .B(n2149), .C(n2148), .ZN(n2150) );
  MUX2ND0 U2586 ( .I0(R_lat_mag[8]), .I1(n2180), .S(n2150), .ZN(
        \mult_x_13/n651 ) );
  NR2D0 U2587 ( .A1(n2155), .A2(n2169), .ZN(n2153) );
  OAI22D0 U2588 ( .A1(n2159), .A2(n2173), .B1(n2151), .B2(n2171), .ZN(n2152)
         );
  AOI211D0 U2589 ( .A1(n2178), .A2(n2250), .B(n2153), .C(n2152), .ZN(n2154) );
  MUX2ND0 U2590 ( .I0(R_lat_mag[8]), .I1(n2180), .S(n2154), .ZN(
        \mult_x_13/n652 ) );
  NR2D0 U2591 ( .A1(n2159), .A2(n2169), .ZN(n2157) );
  OAI22D0 U2592 ( .A1(n2164), .A2(n2173), .B1(n2155), .B2(n2171), .ZN(n2156)
         );
  AOI211D0 U2593 ( .A1(n2178), .A2(n2254), .B(n2157), .C(n2156), .ZN(n2158) );
  MUX2ND0 U2594 ( .I0(R_lat_mag[8]), .I1(n2180), .S(n2158), .ZN(
        \mult_x_13/n653 ) );
  NR2D0 U2595 ( .A1(n2164), .A2(n2169), .ZN(n2161) );
  OAI22D0 U2596 ( .A1(n2172), .A2(n2173), .B1(n2159), .B2(n2171), .ZN(n2160)
         );
  AOI211D0 U2597 ( .A1(n2178), .A2(n2162), .B(n2161), .C(n2160), .ZN(n2163) );
  MUX2ND0 U2598 ( .I0(R_lat_mag[8]), .I1(n2180), .S(n2163), .ZN(
        \mult_x_13/n654 ) );
  NR2D0 U2599 ( .A1(n2172), .A2(n2169), .ZN(n2166) );
  OAI22D0 U2600 ( .A1(n2170), .A2(n2173), .B1(n2164), .B2(n2171), .ZN(n2165)
         );
  MUX2ND0 U2601 ( .I0(R_lat_mag[8]), .I1(n2180), .S(n2168), .ZN(
        \mult_x_13/n655 ) );
  NR2D0 U2602 ( .A1(n2170), .A2(n2169), .ZN(n2176) );
  OAI22D0 U2603 ( .A1(n2174), .A2(n2173), .B1(n2172), .B2(n2171), .ZN(n2175)
         );
  AOI211D0 U2604 ( .A1(n2178), .A2(n2177), .B(n2176), .C(n2175), .ZN(n2179) );
  MUX2ND0 U2605 ( .I0(R_lat_mag[8]), .I1(n2180), .S(n2179), .ZN(
        \mult_x_13/n656 ) );
  MUX2ND0 U2606 ( .I0(R_lat_mag[5]), .I1(\mult_x_13/n660 ), .S(n2182), .ZN(
        \mult_x_13/n661 ) );
  INVD0 U2607 ( .I(n2257), .ZN(n2186) );
  OAI222D0 U2608 ( .A1(n2188), .A2(n2187), .B1(n2186), .B2(n2185), .C1(n2184), 
        .C2(n2183), .ZN(n2189) );
  MUX2ND0 U2609 ( .I0(\mult_x_13/n660 ), .I1(R_lat_mag[5]), .S(n2189), .ZN(
        \mult_x_13/n662 ) );
  AOI22D0 U2610 ( .A1(inv_Q_mag[22]), .A2(n2258), .B1(inv_Q_mag[21]), .B2(
        n2257), .ZN(n2191) );
  CKND2D0 U2611 ( .A1(n2192), .A2(n2191), .ZN(n2193) );
  MUX2ND0 U2612 ( .I0(\mult_x_13/n660 ), .I1(R_lat_mag[5]), .S(n2193), .ZN(
        \mult_x_13/n663 ) );
  AOI22D0 U2613 ( .A1(inv_Q_mag[19]), .A2(n2256), .B1(n2194), .B2(n2255), .ZN(
        n2196) );
  AOI22D0 U2614 ( .A1(inv_Q_mag[21]), .A2(n2258), .B1(inv_Q_mag[20]), .B2(
        n2257), .ZN(n2195) );
  CKND2D0 U2615 ( .A1(n2196), .A2(n2195), .ZN(n2197) );
  MUX2ND0 U2616 ( .I0(\mult_x_13/n660 ), .I1(R_lat_mag[5]), .S(n2197), .ZN(
        \mult_x_13/n664 ) );
  AOI22D0 U2617 ( .A1(inv_Q_mag[18]), .A2(n2256), .B1(n2198), .B2(n2255), .ZN(
        n2200) );
  AOI22D0 U2618 ( .A1(inv_Q_mag[20]), .A2(n2258), .B1(inv_Q_mag[19]), .B2(
        n2257), .ZN(n2199) );
  CKND2D0 U2619 ( .A1(n2200), .A2(n2199), .ZN(n2201) );
  MUX2ND0 U2620 ( .I0(\mult_x_13/n660 ), .I1(R_lat_mag[5]), .S(n2201), .ZN(
        \mult_x_13/n665 ) );
  AOI22D0 U2621 ( .A1(inv_Q_mag[17]), .A2(n2256), .B1(n2202), .B2(n2255), .ZN(
        n2204) );
  AOI22D0 U2622 ( .A1(inv_Q_mag[19]), .A2(n2258), .B1(inv_Q_mag[18]), .B2(
        n2257), .ZN(n2203) );
  MUX2ND0 U2623 ( .I0(\mult_x_13/n660 ), .I1(R_lat_mag[5]), .S(n2205), .ZN(
        \mult_x_13/n666 ) );
  AOI22D0 U2624 ( .A1(inv_Q_mag[16]), .A2(n2256), .B1(n2206), .B2(n2255), .ZN(
        n2208) );
  AOI22D0 U2625 ( .A1(inv_Q_mag[18]), .A2(n2258), .B1(inv_Q_mag[17]), .B2(
        n2257), .ZN(n2207) );
  CKND2D0 U2626 ( .A1(n2208), .A2(n2207), .ZN(n2209) );
  MUX2ND0 U2627 ( .I0(\mult_x_13/n660 ), .I1(R_lat_mag[5]), .S(n2209), .ZN(
        \mult_x_13/n667 ) );
  AOI22D0 U2628 ( .A1(inv_Q_mag[15]), .A2(n2256), .B1(n2210), .B2(n2255), .ZN(
        n2212) );
  AOI22D0 U2629 ( .A1(inv_Q_mag[17]), .A2(n2258), .B1(inv_Q_mag[16]), .B2(
        n2257), .ZN(n2211) );
  CKND2D0 U2630 ( .A1(n2212), .A2(n2211), .ZN(n2213) );
  MUX2ND0 U2631 ( .I0(\mult_x_13/n660 ), .I1(R_lat_mag[5]), .S(n2213), .ZN(
        \mult_x_13/n668 ) );
  AOI22D0 U2632 ( .A1(inv_Q_mag[14]), .A2(n2256), .B1(n2214), .B2(n2255), .ZN(
        n2216) );
  AOI22D0 U2633 ( .A1(inv_Q_mag[16]), .A2(n2258), .B1(inv_Q_mag[15]), .B2(
        n2257), .ZN(n2215) );
  CKND2D0 U2634 ( .A1(n2216), .A2(n2215), .ZN(n2217) );
  MUX2ND0 U2635 ( .I0(\mult_x_13/n660 ), .I1(R_lat_mag[5]), .S(n2217), .ZN(
        \mult_x_13/n669 ) );
  AOI22D0 U2636 ( .A1(inv_Q_mag[15]), .A2(n2258), .B1(n2218), .B2(n2255), .ZN(
        n2220) );
  CKND2D0 U2637 ( .A1(n2220), .A2(n2219), .ZN(n2221) );
  MUX2ND0 U2638 ( .I0(\mult_x_13/n660 ), .I1(R_lat_mag[5]), .S(n2221), .ZN(
        \mult_x_13/n670 ) );
  AOI22D0 U2639 ( .A1(inv_Q_mag[14]), .A2(n2258), .B1(n2222), .B2(n2255), .ZN(
        n2224) );
  AOI22D0 U2640 ( .A1(inv_Q_mag[13]), .A2(n2257), .B1(inv_Q_mag[12]), .B2(
        n2256), .ZN(n2223) );
  MUX2ND0 U2641 ( .I0(\mult_x_13/n660 ), .I1(R_lat_mag[5]), .S(n2225), .ZN(
        \mult_x_13/n671 ) );
  AOI22D0 U2642 ( .A1(n2256), .A2(inv_Q_mag[11]), .B1(n2255), .B2(n2226), .ZN(
        n2228) );
  AOI22D0 U2643 ( .A1(inv_Q_mag[13]), .A2(n2258), .B1(inv_Q_mag[12]), .B2(
        n2257), .ZN(n2227) );
  CKND2D0 U2644 ( .A1(n2228), .A2(n2227), .ZN(n2229) );
  MUX2ND0 U2645 ( .I0(\mult_x_13/n660 ), .I1(R_lat_mag[5]), .S(n2229), .ZN(
        \mult_x_13/n672 ) );
  AOI22D0 U2646 ( .A1(n2256), .A2(inv_Q_mag[10]), .B1(n2255), .B2(n2230), .ZN(
        n2232) );
  AOI22D0 U2647 ( .A1(inv_Q_mag[12]), .A2(n2258), .B1(n2257), .B2(
        inv_Q_mag[11]), .ZN(n2231) );
  CKND2D0 U2648 ( .A1(n2232), .A2(n2231), .ZN(n2233) );
  MUX2ND0 U2649 ( .I0(\mult_x_13/n660 ), .I1(R_lat_mag[5]), .S(n2233), .ZN(
        \mult_x_13/n673 ) );
  AOI22D0 U2650 ( .A1(n2256), .A2(inv_Q_mag[9]), .B1(n2255), .B2(n2234), .ZN(
        n2236) );
  AOI22D0 U2651 ( .A1(n2258), .A2(inv_Q_mag[11]), .B1(n2257), .B2(
        inv_Q_mag[10]), .ZN(n2235) );
  CKND2D0 U2652 ( .A1(n2236), .A2(n2235), .ZN(n2237) );
  MUX2ND0 U2653 ( .I0(\mult_x_13/n660 ), .I1(R_lat_mag[5]), .S(n2237), .ZN(
        \mult_x_13/n674 ) );
  AOI22D0 U2654 ( .A1(n2256), .A2(inv_Q_mag[8]), .B1(n2255), .B2(n2238), .ZN(
        n2240) );
  AOI22D0 U2655 ( .A1(n2258), .A2(inv_Q_mag[10]), .B1(n2257), .B2(inv_Q_mag[9]), .ZN(n2239) );
  CKND2D0 U2656 ( .A1(n2240), .A2(n2239), .ZN(n2241) );
  MUX2ND0 U2657 ( .I0(\mult_x_13/n660 ), .I1(R_lat_mag[5]), .S(n2241), .ZN(
        \mult_x_13/n675 ) );
  AOI22D0 U2658 ( .A1(n2256), .A2(inv_Q_mag[7]), .B1(n2255), .B2(n2242), .ZN(
        n2244) );
  AOI22D0 U2659 ( .A1(n2258), .A2(inv_Q_mag[9]), .B1(n2257), .B2(inv_Q_mag[8]), 
        .ZN(n2243) );
  CKND2D0 U2660 ( .A1(n2244), .A2(n2243), .ZN(n2245) );
  MUX2ND0 U2661 ( .I0(\mult_x_13/n660 ), .I1(R_lat_mag[5]), .S(n2245), .ZN(
        \mult_x_13/n676 ) );
  AOI22D0 U2662 ( .A1(n2256), .A2(inv_Q_mag[6]), .B1(n2255), .B2(n2246), .ZN(
        n2248) );
  AOI22D0 U2663 ( .A1(n2258), .A2(inv_Q_mag[8]), .B1(n2257), .B2(inv_Q_mag[7]), 
        .ZN(n2247) );
  CKND2D0 U2664 ( .A1(n2248), .A2(n2247), .ZN(n2249) );
  MUX2ND0 U2665 ( .I0(\mult_x_13/n660 ), .I1(R_lat_mag[5]), .S(n2249), .ZN(
        \mult_x_13/n677 ) );
  AOI22D0 U2666 ( .A1(n2256), .A2(inv_Q_mag[5]), .B1(n2255), .B2(n2250), .ZN(
        n2252) );
  AOI22D0 U2667 ( .A1(n2258), .A2(inv_Q_mag[7]), .B1(n2257), .B2(inv_Q_mag[6]), 
        .ZN(n2251) );
  CKND2D0 U2668 ( .A1(n2252), .A2(n2251), .ZN(n2253) );
  MUX2ND0 U2669 ( .I0(\mult_x_13/n660 ), .I1(R_lat_mag[5]), .S(n2253), .ZN(
        \mult_x_13/n678 ) );
  AOI22D0 U2670 ( .A1(n2258), .A2(inv_Q_mag[6]), .B1(n2257), .B2(inv_Q_mag[5]), 
        .ZN(n2259) );
  CKND2D0 U2671 ( .A1(n2260), .A2(n2259), .ZN(n2261) );
  MUX2ND0 U2672 ( .I0(\mult_x_13/n660 ), .I1(R_lat_mag[5]), .S(n2261), .ZN(
        \mult_x_13/n679 ) );
  MUX2ND0 U2673 ( .I0(add_tc[23]), .I1(n2263), .S(n2262), .ZN(N97) );
  INVD0 U2674 ( .I(sub_tc[23]), .ZN(n2265) );
  MUX2ND0 U2675 ( .I0(sub_tc[23]), .I1(n2265), .S(n2264), .ZN(N148) );
  INR3D0 U2676 ( .A1(inv_rdy), .B1(state[1]), .B2(n2266), .ZN(next_state[1])
         );
  ND4D0 U2677 ( .A1(n74), .A2(n59), .A3(n58), .A4(n57), .ZN(result_comb[5]) );
  ND4D0 U2678 ( .A1(n74), .A2(n50), .A3(n49), .A4(n48), .ZN(result_comb[8]) );
  ND4D0 U2679 ( .A1(n74), .A2(n47), .A3(n46), .A4(n45), .ZN(result_comb[9]) );
  ND4D0 U2680 ( .A1(n74), .A2(n44), .A3(n43), .A4(n42), .ZN(result_comb[10])
         );
  ND4D0 U2681 ( .A1(n74), .A2(n41), .A3(n40), .A4(n39), .ZN(result_comb[11])
         );
  ND4D0 U2682 ( .A1(n74), .A2(n35), .A3(n34), .A4(n33), .ZN(result_comb[13])
         );
  ND4D0 U2683 ( .A1(n74), .A2(n29), .A3(n28), .A4(n27), .ZN(result_comb[15])
         );
  ND4D0 U2684 ( .A1(n74), .A2(n17), .A3(n16), .A4(n15), .ZN(result_comb[19])
         );
  CMPE42D1 U2685 ( .A(\mult_x_13/n297 ), .B(\mult_x_13/n289 ), .C(
        \mult_x_13/n640 ), .CIX(\mult_x_13/n663 ), .D(\mult_x_13/n293 ), .CO(
        \mult_x_13/n285 ), .COX(\mult_x_13/n284 ), .S(\mult_x_13/n286 ) );
  CMPE42D1 U2686 ( .A(\mult_x_13/n236 ), .B(\mult_x_13/n243 ), .C(
        \mult_x_13/n588 ), .CIX(\mult_x_13/n611 ), .D(\mult_x_13/n239 ), .CO(
        \mult_x_13/n232 ), .COX(\mult_x_13/n231 ), .S(\mult_x_13/n233 ) );
  CMPE42D1 U2687 ( .A(\mult_x_13/n615 ), .B(\mult_x_13/n271 ), .C(
        \mult_x_13/n275 ), .CIX(\mult_x_13/n661 ), .D(\mult_x_13/n638 ), .CO(
        \mult_x_13/n267 ), .COX(\mult_x_13/n266 ), .S(\mult_x_13/n268 ) );
  CMPE42D1 U2688 ( .A(\mult_x_13/n563 ), .B(\mult_x_13/n221 ), .C(
        \mult_x_13/n224 ), .CIX(\mult_x_13/n609 ), .D(\mult_x_13/n586 ), .CO(
        \mult_x_13/n217 ), .COX(\mult_x_13/n216 ), .S(\mult_x_13/n218 ) );
  CMPE42D1 U2689 ( .A(\mult_x_13/n214 ), .B(\mult_x_13/n209 ), .C(
        \mult_x_13/n561 ), .CIX(\mult_x_13/n584 ), .D(\mult_x_13/n211 ), .CO(
        \mult_x_13/n206 ), .COX(\mult_x_13/n205 ), .S(\mult_x_13/n207 ) );
  CMPE42D1 U2690 ( .A(\mult_x_13/n262 ), .B(\mult_x_13/n254 ), .C(
        \mult_x_13/n613 ), .CIX(\mult_x_13/n636 ), .D(\mult_x_13/n258 ), .CO(
        \mult_x_13/n250 ), .COX(\mult_x_13/n249 ), .S(\mult_x_13/n251 ) );
  CMPE42D1 U2691 ( .A(\mult_x_9/n608 ), .B(\mult_x_9/n222 ), .C(
        \mult_x_9/n517 ), .CIX(\mult_x_9/n539 ), .D(\mult_x_9/n219 ), .CO(
        \mult_x_9/n214 ), .COX(\mult_x_9/n203 ), .S(\mult_x_9/n215 ) );
  CMPE42D1 U2692 ( .A(\mult_x_9/n660 ), .B(\mult_x_9/n686 ), .C(
        \mult_x_9/n522 ), .CIX(\mult_x_9/n545 ), .D(\mult_x_9/n272 ), .CO(
        \mult_x_9/n264 ), .COX(\mult_x_9/n247 ), .S(\mult_x_9/n265 ) );
  CMPE42D1 U2693 ( .A(\mult_x_13/n238 ), .B(\mult_x_13/n245 ), .C(
        \mult_x_13/n542 ), .CIX(\mult_x_13/n565 ), .D(\mult_x_13/n242 ), .CO(
        \mult_x_13/n235 ), .COX(\mult_x_13/n234 ), .S(\mult_x_13/n236 ) );
  CMPE42D1 U2694 ( .A(\mult_x_9/n265 ), .B(\mult_x_9/n273 ), .C(
        \mult_x_9/n568 ), .CIX(\mult_x_9/n591 ), .D(\mult_x_9/n269 ), .CO(
        \mult_x_9/n262 ), .COX(\mult_x_9/n261 ), .S(\mult_x_9/n263 ) );
  CMPE42D1 U2695 ( .A(\mult_x_9/n238 ), .B(\mult_x_9/n245 ), .C(
        \mult_x_9/n542 ), .CIX(\mult_x_9/n565 ), .D(\mult_x_9/n242 ), .CO(
        \mult_x_9/n235 ), .COX(\mult_x_9/n234 ), .S(\mult_x_9/n236 ) );
  CMPE42D1 U2696 ( .A(\mult_x_13/n265 ), .B(\mult_x_13/n273 ), .C(
        \mult_x_13/n568 ), .CIX(\mult_x_13/n591 ), .D(\mult_x_13/n269 ), .CO(
        \mult_x_13/n262 ), .COX(\mult_x_13/n261 ), .S(\mult_x_13/n263 ) );
  CMPE42D1 U2697 ( .A(\mult_x_13/n608 ), .B(\mult_x_13/n222 ), .C(
        \mult_x_13/n517 ), .CIX(\mult_x_13/n539 ), .D(\mult_x_13/n219 ), .CO(
        \mult_x_13/n214 ), .COX(\mult_x_13/n203 ), .S(\mult_x_13/n215 ) );
  CMPE42D1 U2698 ( .A(\mult_x_13/n660 ), .B(\mult_x_13/n686 ), .C(
        \mult_x_13/n522 ), .CIX(\mult_x_13/n545 ), .D(\mult_x_13/n272 ), .CO(
        \mult_x_13/n264 ), .COX(\mult_x_13/n247 ), .S(\mult_x_13/n265 ) );
  CMPE42D1 U2699 ( .A(\mult_x_9/n526 ), .B(\mult_x_9/n549 ), .C(
        \mult_x_9/n308 ), .CIX(\mult_x_9/n309 ), .D(\mult_x_9/n572 ), .CO(
        \mult_x_9/n300 ), .COX(\mult_x_9/n299 ), .S(\mult_x_9/n301 ) );
  CMPE42D1 U2700 ( .A(\mult_x_13/n526 ), .B(\mult_x_13/n549 ), .C(
        \mult_x_13/n308 ), .CIX(\mult_x_13/n309 ), .D(\mult_x_13/n572 ), .CO(
        \mult_x_13/n300 ), .COX(\mult_x_13/n299 ), .S(\mult_x_13/n301 ) );
  CMPE42D1 U2701 ( .A(\mult_x_9/n301 ), .B(\mult_x_9/n595 ), .C(
        \mult_x_9/n305 ), .CIX(\mult_x_9/n306 ), .D(\mult_x_9/n618 ), .CO(
        \mult_x_9/n297 ), .COX(\mult_x_9/n296 ), .S(\mult_x_9/n298 ) );
  CMPE42D1 U2702 ( .A(\mult_x_13/n301 ), .B(\mult_x_13/n595 ), .C(
        \mult_x_13/n305 ), .CIX(\mult_x_13/n306 ), .D(\mult_x_13/n618 ), .CO(
        \mult_x_13/n297 ), .COX(\mult_x_13/n296 ), .S(\mult_x_13/n298 ) );
  CMPE42D1 U2703 ( .A(\mult_x_13/n513 ), .B(\mult_x_13/n193 ), .C(
        \mult_x_13/n535 ), .CIX(\mult_x_13/n558 ), .D(\mult_x_13/n194 ), .CO(
        \mult_x_13/n191 ), .COX(\mult_x_13/n190 ), .S(\mult_x_13/n192 ) );
  CMPE42D1 U2704 ( .A(\mult_x_13/n537 ), .B(\mult_x_13/n202 ), .C(
        \mult_x_13/n205 ), .CIX(\mult_x_13/n583 ), .D(\mult_x_13/n560 ), .CO(
        \mult_x_13/n199 ), .COX(\mult_x_13/n198 ), .S(\mult_x_13/n200 ) );
  CMPE42D1 U2705 ( .A(\mult_x_13/n193 ), .B(\mult_x_13/n512 ), .C(
        \mult_x_13/n190 ), .CIX(\mult_x_13/n557 ), .D(\mult_x_13/n534 ), .CO(
        \mult_x_13/n186 ), .COX(\mult_x_13/n185 ), .S(\mult_x_13/n187 ) );
  CMPE42D1 U2706 ( .A(R[2]), .B(\mult_x_9/n523 ), .C(\mult_x_9/n281 ), .CIX(
        \mult_x_9/n282 ), .D(\mult_x_9/n546 ), .CO(\mult_x_9/n273 ), .COX(
        \mult_x_9/n272 ), .S(\mult_x_9/n274 ) );
  CMPE42D1 U2707 ( .A(R_lat_mag[2]), .B(\mult_x_13/n523 ), .C(\mult_x_13/n281 ), .CIX(\mult_x_13/n282 ), .D(\mult_x_13/n546 ), .CO(\mult_x_13/n273 ), .COX(
        \mult_x_13/n272 ), .S(\mult_x_13/n274 ) );
  CMPE42D1 U2708 ( .A(\mult_x_9/n255 ), .B(\mult_x_9/n246 ), .C(
        \mult_x_9/n252 ), .CIX(\mult_x_9/n253 ), .D(\mult_x_9/n566 ), .CO(
        \mult_x_9/n243 ), .COX(\mult_x_9/n242 ), .S(\mult_x_9/n244 ) );
  CMPE42D1 U2709 ( .A(\mult_x_9/n569 ), .B(\mult_x_9/n274 ), .C(
        \mult_x_9/n278 ), .CIX(\mult_x_9/n279 ), .D(\mult_x_9/n592 ), .CO(
        \mult_x_9/n270 ), .COX(\mult_x_9/n269 ), .S(\mult_x_9/n271 ) );
  CMPE42D1 U2710 ( .A(\mult_x_9/n230 ), .B(\mult_x_9/n518 ), .C(
        \mult_x_9/n227 ), .CIX(\mult_x_9/n228 ), .D(\mult_x_9/n540 ), .CO(
        \mult_x_9/n220 ), .COX(\mult_x_9/n219 ), .S(\mult_x_9/n221 ) );
  CMPE42D1 U2711 ( .A(\mult_x_13/n569 ), .B(\mult_x_13/n274 ), .C(
        \mult_x_13/n278 ), .CIX(\mult_x_13/n279 ), .D(\mult_x_13/n592 ), .CO(
        \mult_x_13/n270 ), .COX(\mult_x_13/n269 ), .S(\mult_x_13/n271 ) );
  CMPE42D1 U2712 ( .A(\mult_x_13/n255 ), .B(\mult_x_13/n246 ), .C(
        \mult_x_13/n252 ), .CIX(\mult_x_13/n253 ), .D(\mult_x_13/n566 ), .CO(
        \mult_x_13/n243 ), .COX(\mult_x_13/n242 ), .S(\mult_x_13/n244 ) );
  CMPE42D1 U2713 ( .A(\mult_x_13/n230 ), .B(\mult_x_13/n518 ), .C(
        \mult_x_13/n227 ), .CIX(\mult_x_13/n228 ), .D(\mult_x_13/n540 ), .CO(
        \mult_x_13/n220 ), .COX(\mult_x_13/n219 ), .S(\mult_x_13/n221 ) );
  CMPE42D1 U2714 ( .A(\mult_x_13/n589 ), .B(\mult_x_13/n244 ), .C(
        \mult_x_13/n249 ), .CIX(\mult_x_13/n635 ), .D(\mult_x_13/n612 ), .CO(
        \mult_x_13/n240 ), .COX(\mult_x_13/n239 ), .S(\mult_x_13/n241 ) );
  CMPE42D1 U2715 ( .A(\mult_x_13/n215 ), .B(\mult_x_13/n220 ), .C(
        \mult_x_13/n562 ), .CIX(\mult_x_13/n585 ), .D(\mult_x_13/n216 ), .CO(
        \mult_x_13/n212 ), .COX(\mult_x_13/n211 ), .S(\mult_x_13/n213 ) );
  CMPE42D1 U2716 ( .A(\mult_x_13/n263 ), .B(\mult_x_13/n270 ), .C(
        \mult_x_13/n614 ), .CIX(\mult_x_13/n637 ), .D(\mult_x_13/n266 ), .CO(
        \mult_x_13/n259 ), .COX(\mult_x_13/n258 ), .S(\mult_x_13/n260 ) );
  CMPE42D1 U2717 ( .A(\mult_x_13/n556 ), .B(\mult_x_13/n188 ), .C(
        \mult_x_13/n511 ), .CIX(\mult_x_13/n533 ), .D(\mult_x_13/n185 ), .CO(
        \mult_x_13/n183 ), .COX(\mult_x_13/n178 ), .S(\mult_x_13/n184 ) );
  CMPE42D1 U2718 ( .A(\mult_x_13/n298 ), .B(\mult_x_13/n641 ), .C(
        \mult_x_13/n302 ), .CIX(\mult_x_13/n303 ), .D(\mult_x_13/n664 ), .CO(
        \mult_x_13/n294 ), .COX(\mult_x_13/n293 ), .S(\mult_x_13/n295 ) );
  CMPE42D1 U2719 ( .A(\mult_x_13/n616 ), .B(\mult_x_13/n280 ), .C(
        \mult_x_13/n284 ), .CIX(\mult_x_13/n662 ), .D(\mult_x_13/n639 ), .CO(
        \mult_x_13/n276 ), .COX(\mult_x_13/n275 ), .S(\mult_x_13/n277 ) );
  CMPE42D1 U2720 ( .A(\mult_x_13/n235 ), .B(\mult_x_13/n229 ), .C(
        \mult_x_13/n587 ), .CIX(\mult_x_13/n610 ), .D(\mult_x_13/n231 ), .CO(
        \mult_x_13/n225 ), .COX(\mult_x_13/n224 ), .S(\mult_x_13/n226 ) );
  CMPE42D1 U2721 ( .A(R_lat_mag[2]), .B(\mult_x_13/n525 ), .C(\mult_x_13/n548 ), .CIX(\mult_x_13/n571 ), .D(\mult_x_13/n299 ), .CO(\mult_x_13/n291 ), .COX(
        \mult_x_13/n290 ), .S(\mult_x_13/n292 ) );
  CMPE42D1 U2722 ( .A(\mult_x_13/n300 ), .B(\mult_x_13/n292 ), .C(
        \mult_x_13/n594 ), .CIX(\mult_x_13/n617 ), .D(\mult_x_13/n296 ), .CO(
        \mult_x_13/n288 ), .COX(\mult_x_13/n287 ), .S(\mult_x_13/n289 ) );
  CMPE42D1 U2723 ( .A(\mult_x_13/n237 ), .B(\mult_x_13/n230 ), .C(
        \mult_x_13/n541 ), .CIX(\mult_x_13/n564 ), .D(\mult_x_13/n234 ), .CO(
        \mult_x_13/n228 ), .COX(\mult_x_13/n227 ), .S(\mult_x_13/n229 ) );
  CMPE42D1 U2724 ( .A(\mult_x_9/n264 ), .B(\mult_x_9/n256 ), .C(
        \mult_x_9/n567 ), .CIX(\mult_x_9/n590 ), .D(\mult_x_9/n261 ), .CO(
        \mult_x_9/n253 ), .COX(\mult_x_9/n252 ), .S(\mult_x_9/n254 ) );
  CMPE42D1 U2725 ( .A(R[2]), .B(\mult_x_9/n525 ), .C(\mult_x_9/n548 ), .CIX(
        \mult_x_9/n571 ), .D(\mult_x_9/n299 ), .CO(\mult_x_9/n291 ), .COX(
        \mult_x_9/n290 ), .S(\mult_x_9/n292 ) );
  CMPE42D1 U2726 ( .A(\mult_x_9/n300 ), .B(\mult_x_9/n292 ), .C(
        \mult_x_9/n594 ), .CIX(\mult_x_9/n617 ), .D(\mult_x_9/n296 ), .CO(
        \mult_x_9/n288 ), .COX(\mult_x_9/n287 ), .S(\mult_x_9/n289 ) );
  CMPE42D1 U2727 ( .A(\mult_x_9/n237 ), .B(\mult_x_9/n230 ), .C(
        \mult_x_9/n541 ), .CIX(\mult_x_9/n564 ), .D(\mult_x_9/n234 ), .CO(
        \mult_x_9/n228 ), .COX(\mult_x_9/n227 ), .S(\mult_x_9/n229 ) );
  CMPE42D1 U2728 ( .A(\mult_x_13/n264 ), .B(\mult_x_13/n256 ), .C(
        \mult_x_13/n567 ), .CIX(\mult_x_13/n590 ), .D(\mult_x_13/n261 ), .CO(
        \mult_x_13/n253 ), .COX(\mult_x_13/n252 ), .S(\mult_x_13/n254 ) );
  CMPE42D1 U2729 ( .A(\mult_x_9/n374 ), .B(\mult_x_9/n603 ), .C(
        \mult_x_9/n378 ), .CIX(\mult_x_9/n379 ), .D(\mult_x_9/n626 ), .CO(
        \mult_x_9/n371 ), .COX(\mult_x_9/n370 ), .S(\mult_x_9/n372 ) );
  CMPE42D1 U2730 ( .A(\mult_x_13/n374 ), .B(\mult_x_13/n603 ), .C(
        \mult_x_13/n378 ), .CIX(\mult_x_13/n379 ), .D(\mult_x_13/n626 ), .CO(
        \mult_x_13/n371 ), .COX(\mult_x_13/n370 ), .S(\mult_x_13/n372 ) );
  CMPE42D1 U2731 ( .A(\mult_x_9/n366 ), .B(\mult_x_9/n602 ), .C(
        \mult_x_9/n370 ), .CIX(\mult_x_9/n371 ), .D(\mult_x_9/n625 ), .CO(
        \mult_x_9/n363 ), .COX(\mult_x_9/n362 ), .S(\mult_x_9/n364 ) );
  CMPE42D1 U2732 ( .A(\mult_x_13/n366 ), .B(\mult_x_13/n602 ), .C(
        \mult_x_13/n370 ), .CIX(\mult_x_13/n371 ), .D(\mult_x_13/n625 ), .CO(
        \mult_x_13/n363 ), .COX(\mult_x_13/n362 ), .S(\mult_x_13/n364 ) );
  CMPE42D1 U2733 ( .A(\mult_x_9/n528 ), .B(\mult_x_9/n551 ), .C(
        \mult_x_9/n326 ), .CIX(\mult_x_9/n327 ), .D(\mult_x_9/n574 ), .CO(
        \mult_x_9/n318 ), .COX(\mult_x_9/n317 ), .S(\mult_x_9/n319 ) );
  CMPE42D1 U2734 ( .A(\mult_x_9/n356 ), .B(\mult_x_9/n601 ), .C(
        \mult_x_9/n362 ), .CIX(\mult_x_9/n363 ), .D(\mult_x_9/n624 ), .CO(
        \mult_x_9/n353 ), .COX(\mult_x_9/n352 ), .S(\mult_x_9/n354 ) );
  CMPE42D1 U2735 ( .A(\mult_x_13/n356 ), .B(\mult_x_13/n601 ), .C(
        \mult_x_13/n362 ), .CIX(\mult_x_13/n363 ), .D(\mult_x_13/n624 ), .CO(
        \mult_x_13/n353 ), .COX(\mult_x_13/n352 ), .S(\mult_x_13/n354 ) );
  CMPE42D1 U2736 ( .A(\mult_x_13/n528 ), .B(\mult_x_13/n551 ), .C(
        \mult_x_13/n326 ), .CIX(\mult_x_13/n327 ), .D(\mult_x_13/n574 ), .CO(
        \mult_x_13/n318 ), .COX(\mult_x_13/n317 ), .S(\mult_x_13/n319 ) );
  CMPE42D1 U2737 ( .A(\mult_x_9/n527 ), .B(\mult_x_9/n550 ), .C(
        \mult_x_9/n317 ), .CIX(\mult_x_9/n318 ), .D(\mult_x_9/n573 ), .CO(
        \mult_x_9/n309 ), .COX(\mult_x_9/n308 ), .S(\mult_x_9/n310 ) );
  CMPE42D1 U2738 ( .A(\mult_x_9/n346 ), .B(\mult_x_9/n600 ), .C(
        \mult_x_9/n352 ), .CIX(\mult_x_9/n353 ), .D(\mult_x_9/n623 ), .CO(
        \mult_x_9/n343 ), .COX(\mult_x_9/n342 ), .S(\mult_x_9/n344 ) );
  CMPE42D1 U2739 ( .A(\mult_x_13/n346 ), .B(\mult_x_13/n600 ), .C(
        \mult_x_13/n352 ), .CIX(\mult_x_13/n353 ), .D(\mult_x_13/n623 ), .CO(
        \mult_x_13/n343 ), .COX(\mult_x_13/n342 ), .S(\mult_x_13/n344 ) );
  CMPE42D1 U2740 ( .A(\mult_x_13/n527 ), .B(\mult_x_13/n550 ), .C(
        \mult_x_13/n317 ), .CIX(\mult_x_13/n318 ), .D(\mult_x_13/n573 ), .CO(
        \mult_x_13/n309 ), .COX(\mult_x_13/n308 ), .S(\mult_x_13/n310 ) );
  CMPE42D1 U2741 ( .A(\mult_x_9/n336 ), .B(\mult_x_9/n599 ), .C(
        \mult_x_9/n342 ), .CIX(\mult_x_9/n343 ), .D(\mult_x_9/n622 ), .CO(
        \mult_x_9/n333 ), .COX(\mult_x_9/n332 ), .S(\mult_x_9/n334 ) );
  CMPE42D1 U2742 ( .A(\mult_x_13/n336 ), .B(\mult_x_13/n599 ), .C(
        \mult_x_13/n342 ), .CIX(\mult_x_13/n343 ), .D(\mult_x_13/n622 ), .CO(
        \mult_x_13/n333 ), .COX(\mult_x_13/n332 ), .S(\mult_x_13/n334 ) );
  CMPE42D1 U2743 ( .A(\mult_x_9/n328 ), .B(\mult_x_9/n598 ), .C(
        \mult_x_9/n332 ), .CIX(\mult_x_9/n333 ), .D(\mult_x_9/n621 ), .CO(
        \mult_x_9/n324 ), .COX(\mult_x_9/n323 ), .S(\mult_x_9/n325 ) );
  CMPE42D1 U2744 ( .A(\mult_x_13/n328 ), .B(\mult_x_13/n598 ), .C(
        \mult_x_13/n332 ), .CIX(\mult_x_13/n333 ), .D(\mult_x_13/n621 ), .CO(
        \mult_x_13/n324 ), .COX(\mult_x_13/n323 ), .S(\mult_x_13/n325 ) );
  CMPE42D1 U2745 ( .A(R[2]), .B(\mult_x_9/n524 ), .C(\mult_x_9/n290 ), .CIX(
        \mult_x_9/n291 ), .D(\mult_x_9/n547 ), .CO(\mult_x_9/n282 ), .COX(
        \mult_x_9/n281 ), .S(\mult_x_9/n283 ) );
  CMPE42D1 U2746 ( .A(\mult_x_9/n319 ), .B(\mult_x_9/n597 ), .C(
        \mult_x_9/n323 ), .CIX(\mult_x_9/n324 ), .D(\mult_x_9/n620 ), .CO(
        \mult_x_9/n315 ), .COX(\mult_x_9/n314 ), .S(\mult_x_9/n316 ) );
  CMPE42D1 U2747 ( .A(\mult_x_13/n319 ), .B(\mult_x_13/n597 ), .C(
        \mult_x_13/n323 ), .CIX(\mult_x_13/n324 ), .D(\mult_x_13/n620 ), .CO(
        \mult_x_13/n315 ), .COX(\mult_x_13/n314 ), .S(\mult_x_13/n316 ) );
  CMPE42D1 U2748 ( .A(R_lat_mag[2]), .B(\mult_x_13/n524 ), .C(\mult_x_13/n290 ), .CIX(\mult_x_13/n291 ), .D(\mult_x_13/n547 ), .CO(\mult_x_13/n282 ), .COX(
        \mult_x_13/n281 ), .S(\mult_x_13/n283 ) );
  CMPE42D1 U2749 ( .A(\mult_x_9/n570 ), .B(\mult_x_9/n283 ), .C(
        \mult_x_9/n287 ), .CIX(\mult_x_9/n288 ), .D(\mult_x_9/n593 ), .CO(
        \mult_x_9/n279 ), .COX(\mult_x_9/n278 ), .S(\mult_x_9/n280 ) );
  CMPE42D1 U2750 ( .A(\mult_x_9/n310 ), .B(\mult_x_9/n596 ), .C(
        \mult_x_9/n314 ), .CIX(\mult_x_9/n315 ), .D(\mult_x_9/n619 ), .CO(
        \mult_x_9/n306 ), .COX(\mult_x_9/n305 ), .S(\mult_x_9/n307 ) );
  CMPE42D1 U2751 ( .A(\mult_x_13/n310 ), .B(\mult_x_13/n596 ), .C(
        \mult_x_13/n314 ), .CIX(\mult_x_13/n315 ), .D(\mult_x_13/n619 ), .CO(
        \mult_x_13/n306 ), .COX(\mult_x_13/n305 ), .S(\mult_x_13/n307 ) );
  CMPE42D1 U2752 ( .A(\mult_x_13/n570 ), .B(\mult_x_13/n283 ), .C(
        \mult_x_13/n287 ), .CIX(\mult_x_13/n288 ), .D(\mult_x_13/n593 ), .CO(
        \mult_x_13/n279 ), .COX(\mult_x_13/n278 ), .S(\mult_x_13/n280 ) );
  CMPE42D1 U2753 ( .A(\mult_x_9/n307 ), .B(\mult_x_9/n642 ), .C(
        \mult_x_9/n311 ), .CIX(\mult_x_9/n312 ), .D(\mult_x_9/n665 ), .CO(
        \mult_x_9/n303 ), .COX(\mult_x_9/n302 ), .S(\mult_x_9/n304 ) );
  CMPE42D1 U2754 ( .A(\mult_x_9/n316 ), .B(\mult_x_9/n643 ), .C(
        \mult_x_9/n320 ), .CIX(\mult_x_9/n321 ), .D(\mult_x_9/n666 ), .CO(
        \mult_x_9/n312 ), .COX(\mult_x_9/n311 ), .S(\mult_x_9/n313 ) );
  CMPE42D1 U2755 ( .A(\mult_x_9/n325 ), .B(\mult_x_9/n644 ), .C(
        \mult_x_9/n329 ), .CIX(\mult_x_9/n330 ), .D(\mult_x_9/n667 ), .CO(
        \mult_x_9/n321 ), .COX(\mult_x_9/n320 ), .S(\mult_x_9/n322 ) );
  CMPE42D1 U2756 ( .A(\mult_x_9/n334 ), .B(\mult_x_9/n645 ), .C(
        \mult_x_9/n339 ), .CIX(\mult_x_9/n340 ), .D(\mult_x_9/n668 ), .CO(
        \mult_x_9/n330 ), .COX(\mult_x_9/n329 ), .S(\mult_x_9/n331 ) );
  CMPE42D1 U2757 ( .A(\mult_x_9/n344 ), .B(\mult_x_9/n646 ), .C(
        \mult_x_9/n349 ), .CIX(\mult_x_9/n350 ), .D(\mult_x_9/n669 ), .CO(
        \mult_x_9/n340 ), .COX(\mult_x_9/n339 ), .S(\mult_x_9/n341 ) );
  CMPE42D1 U2758 ( .A(\mult_x_9/n354 ), .B(\mult_x_9/n647 ), .C(
        \mult_x_9/n359 ), .CIX(\mult_x_9/n360 ), .D(\mult_x_9/n670 ), .CO(
        \mult_x_9/n350 ), .COX(\mult_x_9/n349 ), .S(\mult_x_9/n351 ) );
  CMPE42D1 U2759 ( .A(\mult_x_9/n364 ), .B(\mult_x_9/n648 ), .C(
        \mult_x_9/n367 ), .CIX(\mult_x_9/n368 ), .D(\mult_x_9/n671 ), .CO(
        \mult_x_9/n360 ), .COX(\mult_x_9/n359 ), .S(\mult_x_9/n361 ) );
  CMPE42D1 U2760 ( .A(\mult_x_9/n372 ), .B(\mult_x_9/n649 ), .C(
        \mult_x_9/n375 ), .CIX(\mult_x_9/n376 ), .D(\mult_x_9/n672 ), .CO(
        \mult_x_9/n368 ), .COX(\mult_x_9/n367 ), .S(\mult_x_9/n369 ) );
  CMPE42D1 U2761 ( .A(\mult_x_9/n380 ), .B(\mult_x_9/n650 ), .C(
        \mult_x_9/n383 ), .CIX(\mult_x_9/n384 ), .D(\mult_x_9/n673 ), .CO(
        \mult_x_9/n376 ), .COX(\mult_x_9/n375 ), .S(\mult_x_9/n377 ) );
  CMPE42D1 U2762 ( .A(\mult_x_9/n387 ), .B(\mult_x_9/n651 ), .C(
        \mult_x_9/n390 ), .CIX(\mult_x_9/n391 ), .D(\mult_x_9/n674 ), .CO(
        \mult_x_9/n384 ), .COX(\mult_x_9/n383 ), .S(\mult_x_9/n385 ) );
  CMPE42D1 U2763 ( .A(\mult_x_9/n413 ), .B(\mult_x_9/n655 ), .C(
        \mult_x_9/n414 ), .CIX(\mult_x_9/n415 ), .D(\mult_x_9/n678 ), .CO(
        \mult_x_9/n410 ), .COX(\mult_x_9/n409 ), .S(\mult_x_9/n411 ) );
  CMPE42D1 U2764 ( .A(\mult_x_9/n408 ), .B(\mult_x_9/n654 ), .C(
        \mult_x_9/n409 ), .CIX(\mult_x_9/n410 ), .D(\mult_x_9/n677 ), .CO(
        \mult_x_9/n405 ), .COX(\mult_x_9/n404 ), .S(\mult_x_9/n406 ) );
  CMPE42D1 U2765 ( .A(\mult_x_9/n401 ), .B(\mult_x_9/n653 ), .C(
        \mult_x_9/n404 ), .CIX(\mult_x_9/n405 ), .D(\mult_x_9/n676 ), .CO(
        \mult_x_9/n398 ), .COX(\mult_x_9/n397 ), .S(\mult_x_9/n399 ) );
  CMPE42D1 U2766 ( .A(\mult_x_9/n394 ), .B(\mult_x_9/n652 ), .C(
        \mult_x_9/n397 ), .CIX(\mult_x_9/n398 ), .D(\mult_x_9/n675 ), .CO(
        \mult_x_9/n391 ), .COX(\mult_x_9/n390 ), .S(\mult_x_9/n392 ) );
  CMPE42D1 U2767 ( .A(\mult_x_13/n394 ), .B(\mult_x_13/n652 ), .C(
        \mult_x_13/n397 ), .CIX(\mult_x_13/n398 ), .D(\mult_x_13/n675 ), .CO(
        \mult_x_13/n391 ), .COX(\mult_x_13/n390 ), .S(\mult_x_13/n392 ) );
  CMPE42D1 U2768 ( .A(\mult_x_13/n408 ), .B(\mult_x_13/n654 ), .C(
        \mult_x_13/n409 ), .CIX(\mult_x_13/n410 ), .D(\mult_x_13/n677 ), .CO(
        \mult_x_13/n405 ), .COX(\mult_x_13/n404 ), .S(\mult_x_13/n406 ) );
  CMPE42D1 U2769 ( .A(\mult_x_13/n413 ), .B(\mult_x_13/n655 ), .C(
        \mult_x_13/n414 ), .CIX(\mult_x_13/n415 ), .D(\mult_x_13/n678 ), .CO(
        \mult_x_13/n410 ), .COX(\mult_x_13/n409 ), .S(\mult_x_13/n411 ) );
  CMPE42D1 U2770 ( .A(\mult_x_13/n401 ), .B(\mult_x_13/n653 ), .C(
        \mult_x_13/n404 ), .CIX(\mult_x_13/n405 ), .D(\mult_x_13/n676 ), .CO(
        \mult_x_13/n398 ), .COX(\mult_x_13/n397 ), .S(\mult_x_13/n399 ) );
  CMPE42D1 U2771 ( .A(\mult_x_13/n387 ), .B(\mult_x_13/n651 ), .C(
        \mult_x_13/n390 ), .CIX(\mult_x_13/n391 ), .D(\mult_x_13/n674 ), .CO(
        \mult_x_13/n384 ), .COX(\mult_x_13/n383 ), .S(\mult_x_13/n385 ) );
  CMPE42D1 U2772 ( .A(\mult_x_13/n380 ), .B(\mult_x_13/n650 ), .C(
        \mult_x_13/n383 ), .CIX(\mult_x_13/n384 ), .D(\mult_x_13/n673 ), .CO(
        \mult_x_13/n376 ), .COX(\mult_x_13/n375 ), .S(\mult_x_13/n377 ) );
  CMPE42D1 U2773 ( .A(\mult_x_13/n372 ), .B(\mult_x_13/n649 ), .C(
        \mult_x_13/n375 ), .CIX(\mult_x_13/n376 ), .D(\mult_x_13/n672 ), .CO(
        \mult_x_13/n368 ), .COX(\mult_x_13/n367 ), .S(\mult_x_13/n369 ) );
  CMPE42D1 U2774 ( .A(\mult_x_13/n364 ), .B(\mult_x_13/n648 ), .C(
        \mult_x_13/n367 ), .CIX(\mult_x_13/n368 ), .D(\mult_x_13/n671 ), .CO(
        \mult_x_13/n360 ), .COX(\mult_x_13/n359 ), .S(\mult_x_13/n361 ) );
  CMPE42D1 U2775 ( .A(\mult_x_13/n354 ), .B(\mult_x_13/n647 ), .C(
        \mult_x_13/n359 ), .CIX(\mult_x_13/n360 ), .D(\mult_x_13/n670 ), .CO(
        \mult_x_13/n350 ), .COX(\mult_x_13/n349 ), .S(\mult_x_13/n351 ) );
  CMPE42D1 U2776 ( .A(\mult_x_13/n344 ), .B(\mult_x_13/n646 ), .C(
        \mult_x_13/n349 ), .CIX(\mult_x_13/n350 ), .D(\mult_x_13/n669 ), .CO(
        \mult_x_13/n340 ), .COX(\mult_x_13/n339 ), .S(\mult_x_13/n341 ) );
  CMPE42D1 U2777 ( .A(\mult_x_13/n334 ), .B(\mult_x_13/n645 ), .C(
        \mult_x_13/n339 ), .CIX(\mult_x_13/n340 ), .D(\mult_x_13/n668 ), .CO(
        \mult_x_13/n330 ), .COX(\mult_x_13/n329 ), .S(\mult_x_13/n331 ) );
  CMPE42D1 U2778 ( .A(\mult_x_13/n325 ), .B(\mult_x_13/n644 ), .C(
        \mult_x_13/n329 ), .CIX(\mult_x_13/n330 ), .D(\mult_x_13/n667 ), .CO(
        \mult_x_13/n321 ), .COX(\mult_x_13/n320 ), .S(\mult_x_13/n322 ) );
  CMPE42D1 U2779 ( .A(\mult_x_13/n316 ), .B(\mult_x_13/n643 ), .C(
        \mult_x_13/n320 ), .CIX(\mult_x_13/n321 ), .D(\mult_x_13/n666 ), .CO(
        \mult_x_13/n312 ), .COX(\mult_x_13/n311 ), .S(\mult_x_13/n313 ) );
  CMPE42D1 U2780 ( .A(\mult_x_13/n307 ), .B(\mult_x_13/n642 ), .C(
        \mult_x_13/n311 ), .CIX(\mult_x_13/n312 ), .D(\mult_x_13/n665 ), .CO(
        \mult_x_13/n303 ), .COX(\mult_x_13/n302 ), .S(\mult_x_13/n304 ) );
  CMPE42D1 U2781 ( .A(\mult_x_9/n382 ), .B(\mult_x_9/n604 ), .C(
        \mult_x_9/n388 ), .CIX(\mult_x_9/n386 ), .D(\mult_x_9/n627 ), .CO(
        \mult_x_9/n379 ), .COX(\mult_x_9/n378 ), .S(\mult_x_9/n380 ) );
  CMPE42D1 U2782 ( .A(\mult_x_13/n382 ), .B(\mult_x_13/n604 ), .C(
        \mult_x_13/n388 ), .CIX(\mult_x_13/n386 ), .D(\mult_x_13/n627 ), .CO(
        \mult_x_13/n379 ), .COX(\mult_x_13/n378 ), .S(\mult_x_13/n380 ) );
  CMPE42D1 U2783 ( .A(\mult_x_9/n529 ), .B(\mult_x_9/n552 ), .C(
        \mult_x_9/n337 ), .CIX(\mult_x_9/n335 ), .D(\mult_x_9/n575 ), .CO(
        \mult_x_9/n327 ), .COX(\mult_x_9/n326 ), .S(\mult_x_9/n328 ) );
  CMPE42D1 U2784 ( .A(\mult_x_13/n529 ), .B(\mult_x_13/n552 ), .C(
        \mult_x_13/n337 ), .CIX(\mult_x_13/n335 ), .D(\mult_x_13/n575 ), .CO(
        \mult_x_13/n327 ), .COX(\mult_x_13/n326 ), .S(\mult_x_13/n328 ) );
  CMPE42D1 U2785 ( .A(\mult_x_9/n418 ), .B(\mult_x_9/n656 ), .C(
        \mult_x_9/n421 ), .CIX(\mult_x_9/n419 ), .D(\mult_x_9/n679 ), .CO(
        \mult_x_9/n415 ), .COX(\mult_x_9/n414 ), .S(\mult_x_9/n416 ) );
  CMPE42D1 U2786 ( .A(\mult_x_13/n418 ), .B(\mult_x_13/n656 ), .C(
        \mult_x_13/n421 ), .CIX(\mult_x_13/n419 ), .D(\mult_x_13/n679 ), .CO(
        \mult_x_13/n415 ), .COX(\mult_x_13/n414 ), .S(\mult_x_13/n416 ) );
  CMPE42D1 U2787 ( .A(\mult_x_9/n615 ), .B(\mult_x_9/n271 ), .C(
        \mult_x_9/n275 ), .CIX(\mult_x_9/n661 ), .D(\mult_x_9/n638 ), .CO(
        \mult_x_9/n267 ), .COX(\mult_x_9/n266 ), .S(\mult_x_9/n268 ) );
  CMPE42D1 U2788 ( .A(\mult_x_9/n616 ), .B(\mult_x_9/n280 ), .C(
        \mult_x_9/n284 ), .CIX(\mult_x_9/n662 ), .D(\mult_x_9/n639 ), .CO(
        \mult_x_9/n276 ), .COX(\mult_x_9/n275 ), .S(\mult_x_9/n277 ) );
  CMPE42D1 U2789 ( .A(\mult_x_9/n193 ), .B(\mult_x_9/n512 ), .C(
        \mult_x_9/n190 ), .CIX(\mult_x_9/n557 ), .D(\mult_x_9/n534 ), .CO(
        \mult_x_9/n186 ), .COX(\mult_x_9/n185 ), .S(\mult_x_9/n187 ) );
  CMPE42D1 U2790 ( .A(\mult_x_9/n513 ), .B(\mult_x_9/n193 ), .C(
        \mult_x_9/n535 ), .CIX(\mult_x_9/n558 ), .D(\mult_x_9/n194 ), .CO(
        \mult_x_9/n191 ), .COX(\mult_x_9/n190 ), .S(\mult_x_9/n192 ) );
  CMPE42D1 U2791 ( .A(\mult_x_9/n563 ), .B(\mult_x_9/n221 ), .C(
        \mult_x_9/n224 ), .CIX(\mult_x_9/n609 ), .D(\mult_x_9/n586 ), .CO(
        \mult_x_9/n217 ), .COX(\mult_x_9/n216 ), .S(\mult_x_9/n218 ) );
  CMPE42D1 U2792 ( .A(\mult_x_9/n235 ), .B(\mult_x_9/n229 ), .C(
        \mult_x_9/n587 ), .CIX(\mult_x_9/n610 ), .D(\mult_x_9/n231 ), .CO(
        \mult_x_9/n225 ), .COX(\mult_x_9/n224 ), .S(\mult_x_9/n226 ) );
  CMPE42D1 U2793 ( .A(\mult_x_13/n197 ), .B(\mult_x_13/n201 ), .C(
        \mult_x_13/n536 ), .CIX(\mult_x_13/n559 ), .D(\mult_x_13/n198 ), .CO(
        \mult_x_13/n195 ), .COX(\mult_x_13/n194 ), .S(\mult_x_13/n196 ) );
  CMPE42D1 U2794 ( .A(\mult_x_9/n537 ), .B(\mult_x_9/n202 ), .C(
        \mult_x_9/n205 ), .CIX(\mult_x_9/n583 ), .D(\mult_x_9/n560 ), .CO(
        \mult_x_9/n199 ), .COX(\mult_x_9/n198 ), .S(\mult_x_9/n200 ) );
  CMPE42D1 U2795 ( .A(\mult_x_9/n214 ), .B(\mult_x_9/n209 ), .C(
        \mult_x_9/n561 ), .CIX(\mult_x_9/n584 ), .D(\mult_x_9/n211 ), .CO(
        \mult_x_9/n206 ), .COX(\mult_x_9/n205 ), .S(\mult_x_9/n207 ) );
  CMPE42D1 U2796 ( .A(\mult_x_9/n589 ), .B(\mult_x_9/n244 ), .C(
        \mult_x_9/n249 ), .CIX(\mult_x_9/n635 ), .D(\mult_x_9/n612 ), .CO(
        \mult_x_9/n240 ), .COX(\mult_x_9/n239 ), .S(\mult_x_9/n241 ) );
  CMPE42D1 U2797 ( .A(\mult_x_9/n262 ), .B(\mult_x_9/n254 ), .C(
        \mult_x_9/n613 ), .CIX(\mult_x_9/n636 ), .D(\mult_x_9/n258 ), .CO(
        \mult_x_9/n250 ), .COX(\mult_x_9/n249 ), .S(\mult_x_9/n251 ) );
  CMPE42D1 U2798 ( .A(\mult_x_9/n556 ), .B(\mult_x_9/n188 ), .C(
        \mult_x_9/n511 ), .CIX(\mult_x_9/n533 ), .D(\mult_x_9/n185 ), .CO(
        \mult_x_9/n183 ), .COX(\mult_x_9/n178 ), .S(\mult_x_9/n184 ) );
  CMPE42D1 U2799 ( .A(\mult_x_9/n263 ), .B(\mult_x_9/n270 ), .C(
        \mult_x_9/n614 ), .CIX(\mult_x_9/n637 ), .D(\mult_x_9/n266 ), .CO(
        \mult_x_9/n259 ), .COX(\mult_x_9/n258 ), .S(\mult_x_9/n260 ) );
  CMPE42D1 U2800 ( .A(\mult_x_9/n215 ), .B(\mult_x_9/n220 ), .C(
        \mult_x_9/n562 ), .CIX(\mult_x_9/n585 ), .D(\mult_x_9/n216 ), .CO(
        \mult_x_9/n212 ), .COX(\mult_x_9/n211 ), .S(\mult_x_9/n213 ) );
  CMPE42D1 U2801 ( .A(\mult_x_9/n297 ), .B(\mult_x_9/n289 ), .C(
        \mult_x_9/n640 ), .CIX(\mult_x_9/n663 ), .D(\mult_x_9/n293 ), .CO(
        \mult_x_9/n285 ), .COX(\mult_x_9/n284 ), .S(\mult_x_9/n286 ) );
  CMPE42D1 U2802 ( .A(\mult_x_9/n197 ), .B(\mult_x_9/n201 ), .C(
        \mult_x_9/n536 ), .CIX(\mult_x_9/n559 ), .D(\mult_x_9/n198 ), .CO(
        \mult_x_9/n195 ), .COX(\mult_x_9/n194 ), .S(\mult_x_9/n196 ) );
  CMPE42D1 U2803 ( .A(\mult_x_9/n236 ), .B(\mult_x_9/n243 ), .C(
        \mult_x_9/n588 ), .CIX(\mult_x_9/n611 ), .D(\mult_x_9/n239 ), .CO(
        \mult_x_9/n232 ), .COX(\mult_x_9/n231 ), .S(\mult_x_9/n233 ) );
  CMPE42D1 U2804 ( .A(\mult_x_9/n298 ), .B(\mult_x_9/n641 ), .C(
        \mult_x_9/n302 ), .CIX(\mult_x_9/n303 ), .D(\mult_x_9/n664 ), .CO(
        \mult_x_9/n294 ), .COX(\mult_x_9/n293 ), .S(\mult_x_9/n295 ) );
endmodule
