// Created by ihdl
module mult_inv ( clk, rst_n, start, S_mag, Q_mag, rdy );
  input [22:0] S_mag;
  output [22:0] Q_mag;
  input clk, rst_n, start;
  output rdy;
  wire   running, N67, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, \DP_OP_13J3_123_8774/n889 ,
         \DP_OP_13J3_123_8774/n888 , \DP_OP_13J3_123_8774/n887 ,
         \DP_OP_13J3_123_8774/n886 , \DP_OP_13J3_123_8774/n885 ,
         \DP_OP_13J3_123_8774/n884 , \DP_OP_13J3_123_8774/n883 ,
         \DP_OP_13J3_123_8774/n882 , \DP_OP_13J3_123_8774/n881 ,
         \DP_OP_13J3_123_8774/n880 , \DP_OP_13J3_123_8774/n879 ,
         \DP_OP_13J3_123_8774/n878 , \DP_OP_13J3_123_8774/n877 ,
         \DP_OP_13J3_123_8774/n876 , \DP_OP_13J3_123_8774/n875 ,
         \DP_OP_13J3_123_8774/n874 , \DP_OP_13J3_123_8774/n873 ,
         \DP_OP_13J3_123_8774/n872 , \DP_OP_13J3_123_8774/n871 ,
         \DP_OP_13J3_123_8774/n866 , \DP_OP_13J3_123_8774/n865 ,
         \DP_OP_13J3_123_8774/n864 , \DP_OP_13J3_123_8774/n863 ,
         \DP_OP_13J3_123_8774/n862 , \DP_OP_13J3_123_8774/n861 ,
         \DP_OP_13J3_123_8774/n860 , \DP_OP_13J3_123_8774/n859 ,
         \DP_OP_13J3_123_8774/n858 , \DP_OP_13J3_123_8774/n857 ,
         \DP_OP_13J3_123_8774/n856 , \DP_OP_13J3_123_8774/n855 ,
         \DP_OP_13J3_123_8774/n854 , \DP_OP_13J3_123_8774/n853 ,
         \DP_OP_13J3_123_8774/n852 , \DP_OP_13J3_123_8774/n851 ,
         \DP_OP_13J3_123_8774/n850 , \DP_OP_13J3_123_8774/n849 ,
         \DP_OP_13J3_123_8774/n848 , \DP_OP_13J3_123_8774/n847 ,
         \DP_OP_13J3_123_8774/n846 , \DP_OP_13J3_123_8774/n845 ,
         \DP_OP_13J3_123_8774/n837 , \DP_OP_13J3_123_8774/n836 ,
         \DP_OP_13J3_123_8774/n835 , \DP_OP_13J3_123_8774/n834 ,
         \DP_OP_13J3_123_8774/n833 , \DP_OP_13J3_123_8774/n832 ,
         \DP_OP_13J3_123_8774/n831 , \DP_OP_13J3_123_8774/n830 ,
         \DP_OP_13J3_123_8774/n829 , \DP_OP_13J3_123_8774/n828 ,
         \DP_OP_13J3_123_8774/n827 , \DP_OP_13J3_123_8774/n826 ,
         \DP_OP_13J3_123_8774/n825 , \DP_OP_13J3_123_8774/n824 ,
         \DP_OP_13J3_123_8774/n823 , \DP_OP_13J3_123_8774/n822 ,
         \DP_OP_13J3_123_8774/n821 , \DP_OP_13J3_123_8774/n820 ,
         \DP_OP_13J3_123_8774/n819 , \DP_OP_13J3_123_8774/n814 ,
         \DP_OP_13J3_123_8774/n813 , \DP_OP_13J3_123_8774/n812 ,
         \DP_OP_13J3_123_8774/n811 , \DP_OP_13J3_123_8774/n810 ,
         \DP_OP_13J3_123_8774/n809 , \DP_OP_13J3_123_8774/n808 ,
         \DP_OP_13J3_123_8774/n807 , \DP_OP_13J3_123_8774/n806 ,
         \DP_OP_13J3_123_8774/n805 , \DP_OP_13J3_123_8774/n804 ,
         \DP_OP_13J3_123_8774/n803 , \DP_OP_13J3_123_8774/n802 ,
         \DP_OP_13J3_123_8774/n801 , \DP_OP_13J3_123_8774/n800 ,
         \DP_OP_13J3_123_8774/n799 , \DP_OP_13J3_123_8774/n798 ,
         \DP_OP_13J3_123_8774/n797 , \DP_OP_13J3_123_8774/n796 ,
         \DP_OP_13J3_123_8774/n795 , \DP_OP_13J3_123_8774/n794 ,
         \DP_OP_13J3_123_8774/n793 , \DP_OP_13J3_123_8774/n785 ,
         \DP_OP_13J3_123_8774/n784 , \DP_OP_13J3_123_8774/n783 ,
         \DP_OP_13J3_123_8774/n782 , \DP_OP_13J3_123_8774/n781 ,
         \DP_OP_13J3_123_8774/n780 , \DP_OP_13J3_123_8774/n779 ,
         \DP_OP_13J3_123_8774/n778 , \DP_OP_13J3_123_8774/n777 ,
         \DP_OP_13J3_123_8774/n776 , \DP_OP_13J3_123_8774/n775 ,
         \DP_OP_13J3_123_8774/n774 , \DP_OP_13J3_123_8774/n773 ,
         \DP_OP_13J3_123_8774/n772 , \DP_OP_13J3_123_8774/n771 ,
         \DP_OP_13J3_123_8774/n770 , \DP_OP_13J3_123_8774/n769 ,
         \DP_OP_13J3_123_8774/n768 , \DP_OP_13J3_123_8774/n767 ,
         \DP_OP_13J3_123_8774/n762 , \DP_OP_13J3_123_8774/n761 ,
         \DP_OP_13J3_123_8774/n760 , \DP_OP_13J3_123_8774/n759 ,
         \DP_OP_13J3_123_8774/n758 , \DP_OP_13J3_123_8774/n757 ,
         \DP_OP_13J3_123_8774/n756 , \DP_OP_13J3_123_8774/n755 ,
         \DP_OP_13J3_123_8774/n752 , \DP_OP_13J3_123_8774/n751 ,
         \DP_OP_13J3_123_8774/n750 , \DP_OP_13J3_123_8774/n749 ,
         \DP_OP_13J3_123_8774/n747 , \DP_OP_13J3_123_8774/n746 ,
         \DP_OP_13J3_123_8774/n745 , \DP_OP_13J3_123_8774/n744 ,
         \DP_OP_13J3_123_8774/n743 , \DP_OP_13J3_123_8774/n739 ,
         \DP_OP_13J3_123_8774/n738 , \DP_OP_13J3_123_8774/n737 ,
         \DP_OP_13J3_123_8774/n736 , \DP_OP_13J3_123_8774/n735 ,
         \DP_OP_13J3_123_8774/n734 , \DP_OP_13J3_123_8774/n733 ,
         \DP_OP_13J3_123_8774/n732 , \DP_OP_13J3_123_8774/n728 ,
         \DP_OP_13J3_123_8774/n727 , \DP_OP_13J3_123_8774/n723 ,
         \DP_OP_13J3_123_8774/n722 , \DP_OP_13J3_123_8774/n721 ,
         \DP_OP_13J3_123_8774/n631 , \DP_OP_13J3_123_8774/n629 ,
         \DP_OP_13J3_123_8774/n628 , \DP_OP_13J3_123_8774/n626 ,
         \DP_OP_13J3_123_8774/n625 , \DP_OP_13J3_123_8774/n624 ,
         \DP_OP_13J3_123_8774/n623 , \DP_OP_13J3_123_8774/n621 ,
         \DP_OP_13J3_123_8774/n620 , \DP_OP_13J3_123_8774/n619 ,
         \DP_OP_13J3_123_8774/n618 , \DP_OP_13J3_123_8774/n616 ,
         \DP_OP_13J3_123_8774/n615 , \DP_OP_13J3_123_8774/n614 ,
         \DP_OP_13J3_123_8774/n611 , \DP_OP_13J3_123_8774/n609 ,
         \DP_OP_13J3_123_8774/n608 , \DP_OP_13J3_123_8774/n607 ,
         \DP_OP_13J3_123_8774/n604 , \DP_OP_13J3_123_8774/n602 ,
         \DP_OP_13J3_123_8774/n601 , \DP_OP_13J3_123_8774/n600 ,
         \DP_OP_13J3_123_8774/n598 , \DP_OP_13J3_123_8774/n597 ,
         \DP_OP_13J3_123_8774/n596 , \DP_OP_13J3_123_8774/n595 ,
         \DP_OP_13J3_123_8774/n594 , \DP_OP_13J3_123_8774/n593 ,
         \DP_OP_13J3_123_8774/n592 , \DP_OP_13J3_123_8774/n590 ,
         \DP_OP_13J3_123_8774/n589 , \DP_OP_13J3_123_8774/n588 ,
         \DP_OP_13J3_123_8774/n587 , \DP_OP_13J3_123_8774/n586 ,
         \DP_OP_13J3_123_8774/n585 , \DP_OP_13J3_123_8774/n584 ,
         \DP_OP_13J3_123_8774/n582 , \DP_OP_13J3_123_8774/n581 ,
         \DP_OP_13J3_123_8774/n580 , \DP_OP_13J3_123_8774/n579 ,
         \DP_OP_13J3_123_8774/n578 , \DP_OP_13J3_123_8774/n577 ,
         \DP_OP_13J3_123_8774/n576 , \DP_OP_13J3_123_8774/n574 ,
         \DP_OP_13J3_123_8774/n573 , \DP_OP_13J3_123_8774/n572 ,
         \DP_OP_13J3_123_8774/n571 , \DP_OP_13J3_123_8774/n570 ,
         \DP_OP_13J3_123_8774/n569 , \DP_OP_13J3_123_8774/n566 ,
         \DP_OP_13J3_123_8774/n564 , \DP_OP_13J3_123_8774/n563 ,
         \DP_OP_13J3_123_8774/n562 , \DP_OP_13J3_123_8774/n561 ,
         \DP_OP_13J3_123_8774/n560 , \DP_OP_13J3_123_8774/n559 ,
         \DP_OP_13J3_123_8774/n556 , \DP_OP_13J3_123_8774/n554 ,
         \DP_OP_13J3_123_8774/n553 , \DP_OP_13J3_123_8774/n552 ,
         \DP_OP_13J3_123_8774/n551 , \DP_OP_13J3_123_8774/n550 ,
         \DP_OP_13J3_123_8774/n549 , \DP_OP_13J3_123_8774/n547 ,
         \DP_OP_13J3_123_8774/n546 , \DP_OP_13J3_123_8774/n545 ,
         \DP_OP_13J3_123_8774/n544 , \DP_OP_13J3_123_8774/n543 ,
         \DP_OP_13J3_123_8774/n542 , \DP_OP_13J3_123_8774/n541 ,
         \DP_OP_13J3_123_8774/n540 , \DP_OP_13J3_123_8774/n539 ,
         \DP_OP_13J3_123_8774/n538 , \DP_OP_13J3_123_8774/n537 ,
         \DP_OP_13J3_123_8774/n536 , \DP_OP_13J3_123_8774/n535 ,
         \DP_OP_13J3_123_8774/n534 , \DP_OP_13J3_123_8774/n533 ,
         \DP_OP_13J3_123_8774/n532 , \DP_OP_13J3_123_8774/n531 ,
         \DP_OP_13J3_123_8774/n530 , \DP_OP_13J3_123_8774/n529 ,
         \DP_OP_13J3_123_8774/n528 , \DP_OP_13J3_123_8774/n527 ,
         \DP_OP_13J3_123_8774/n526 , \DP_OP_13J3_123_8774/n525 ,
         \DP_OP_13J3_123_8774/n524 , \DP_OP_13J3_123_8774/n523 ,
         \DP_OP_13J3_123_8774/n522 , \DP_OP_13J3_123_8774/n521 ,
         \DP_OP_13J3_123_8774/n520 , \DP_OP_13J3_123_8774/n519 ,
         \DP_OP_13J3_123_8774/n518 , \DP_OP_13J3_123_8774/n517 ,
         \DP_OP_13J3_123_8774/n516 , \DP_OP_13J3_123_8774/n515 ,
         \DP_OP_13J3_123_8774/n514 , \DP_OP_13J3_123_8774/n513 ,
         \DP_OP_13J3_123_8774/n512 , \DP_OP_13J3_123_8774/n511 ,
         \DP_OP_13J3_123_8774/n510 , \DP_OP_13J3_123_8774/n509 ,
         \DP_OP_13J3_123_8774/n508 , \DP_OP_13J3_123_8774/n507 ,
         \DP_OP_13J3_123_8774/n506 , \DP_OP_13J3_123_8774/n505 ,
         \DP_OP_13J3_123_8774/n504 , \DP_OP_13J3_123_8774/n503 ,
         \DP_OP_13J3_123_8774/n502 , \DP_OP_13J3_123_8774/n501 ,
         \DP_OP_13J3_123_8774/n500 , \DP_OP_13J3_123_8774/n499 ,
         \DP_OP_13J3_123_8774/n498 , \DP_OP_13J3_123_8774/n497 ,
         \DP_OP_13J3_123_8774/n496 , \DP_OP_13J3_123_8774/n495 ,
         \DP_OP_13J3_123_8774/n494 , \DP_OP_13J3_123_8774/n493 ,
         \DP_OP_13J3_123_8774/n492 , \DP_OP_13J3_123_8774/n491 ,
         \DP_OP_13J3_123_8774/n490 , \DP_OP_13J3_123_8774/n489 ,
         \DP_OP_13J3_123_8774/n488 , \DP_OP_13J3_123_8774/n487 ,
         \DP_OP_13J3_123_8774/n486 , \DP_OP_13J3_123_8774/n485 ,
         \DP_OP_13J3_123_8774/n484 , \DP_OP_13J3_123_8774/n483 ,
         \DP_OP_13J3_123_8774/n482 , \DP_OP_13J3_123_8774/n481 ,
         \DP_OP_13J3_123_8774/n480 , \DP_OP_13J3_123_8774/n479 ,
         \DP_OP_13J3_123_8774/n478 , \DP_OP_13J3_123_8774/n477 ,
         \DP_OP_13J3_123_8774/n476 , \DP_OP_13J3_123_8774/n475 ,
         \DP_OP_13J3_123_8774/n474 , \DP_OP_13J3_123_8774/n473 ,
         \DP_OP_13J3_123_8774/n472 , \DP_OP_13J3_123_8774/n471 ,
         \DP_OP_13J3_123_8774/n470 , \DP_OP_13J3_123_8774/n469 ,
         \DP_OP_13J3_123_8774/n468 , \DP_OP_13J3_123_8774/n466 ,
         \DP_OP_13J3_123_8774/n465 , \DP_OP_13J3_123_8774/n464 ,
         \DP_OP_13J3_123_8774/n463 , \DP_OP_13J3_123_8774/n462 ,
         \DP_OP_13J3_123_8774/n461 , \DP_OP_13J3_123_8774/n460 ,
         \DP_OP_13J3_123_8774/n459 , \DP_OP_13J3_123_8774/n457 ,
         \DP_OP_13J3_123_8774/n456 , \DP_OP_13J3_123_8774/n455 ,
         \DP_OP_13J3_123_8774/n454 , \DP_OP_13J3_123_8774/n453 ,
         \DP_OP_13J3_123_8774/n452 , \DP_OP_13J3_123_8774/n451 ,
         \DP_OP_13J3_123_8774/n450 , \DP_OP_13J3_123_8774/n449 ,
         \DP_OP_13J3_123_8774/n448 , \DP_OP_13J3_123_8774/n447 ,
         \DP_OP_13J3_123_8774/n446 , \DP_OP_13J3_123_8774/n445 ,
         \DP_OP_13J3_123_8774/n444 , \DP_OP_13J3_123_8774/n443 ,
         \DP_OP_13J3_123_8774/n442 , \DP_OP_13J3_123_8774/n441 ,
         \DP_OP_13J3_123_8774/n440 , \DP_OP_13J3_123_8774/n439 ,
         \DP_OP_13J3_123_8774/n438 , \DP_OP_13J3_123_8774/n437 ,
         \DP_OP_13J3_123_8774/n436 , \DP_OP_13J3_123_8774/n435 ,
         \DP_OP_13J3_123_8774/n434 , \DP_OP_13J3_123_8774/n432 ,
         \DP_OP_13J3_123_8774/n431 , \DP_OP_13J3_123_8774/n430 ,
         \DP_OP_13J3_123_8774/n429 , \DP_OP_13J3_123_8774/n428 ,
         \DP_OP_13J3_123_8774/n427 , \DP_OP_13J3_123_8774/n426 ,
         \DP_OP_13J3_123_8774/n425 , \DP_OP_13J3_123_8774/n424 ,
         \DP_OP_13J3_123_8774/n423 , \DP_OP_13J3_123_8774/n422 ,
         \DP_OP_13J3_123_8774/n421 , \DP_OP_13J3_123_8774/n419 ,
         \DP_OP_13J3_123_8774/n417 , \DP_OP_13J3_123_8774/n416 ,
         \DP_OP_13J3_123_8774/n415 , \DP_OP_13J3_123_8774/n413 ,
         \DP_OP_13J3_123_8774/n412 , \DP_OP_13J3_123_8774/n411 ,
         \DP_OP_13J3_123_8774/n410 , \DP_OP_13J3_123_8774/n409 ,
         \DP_OP_13J3_123_8774/n408 , \DP_OP_13J3_123_8774/n407 ,
         \DP_OP_13J3_123_8774/n406 , \DP_OP_13J3_123_8774/n405 ,
         \DP_OP_13J3_123_8774/n404 , \DP_OP_13J3_123_8774/n403 ,
         \DP_OP_13J3_123_8774/n402 , \DP_OP_13J3_123_8774/n401 ,
         \DP_OP_13J3_123_8774/n400 , \DP_OP_13J3_123_8774/n398 ,
         \DP_OP_13J3_123_8774/n397 , \DP_OP_13J3_123_8774/n396 ,
         \DP_OP_13J3_123_8774/n395 , \DP_OP_13J3_123_8774/n394 ,
         \DP_OP_13J3_123_8774/n393 , \DP_OP_13J3_123_8774/n388 , n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032;
  wire   [4:0] bit_pos;

  DFCNQD1 \bit_pos_reg[0]  ( .D(n74), .CP(clk), .CDN(rst_n), .Q(bit_pos[0]) );
  DFCNQD1 running_reg ( .D(n72), .CP(clk), .CDN(rst_n), .Q(running) );
  DFCNQD1 rdy_reg ( .D(N67), .CP(clk), .CDN(rst_n), .Q(rdy) );
  DFCNQD1 \bit_pos_reg[4]  ( .D(n73), .CP(clk), .CDN(rst_n), .Q(bit_pos[4]) );
  DFCNQD1 \bit_pos_reg[1]  ( .D(n71), .CP(clk), .CDN(rst_n), .Q(bit_pos[1]) );
  DFCNQD1 \bit_pos_reg[2]  ( .D(n70), .CP(clk), .CDN(rst_n), .Q(bit_pos[2]) );
  DFCNQD1 \bit_pos_reg[3]  ( .D(n69), .CP(clk), .CDN(rst_n), .Q(bit_pos[3]) );
  DFCNQD1 \Q_mag_reg[9]  ( .D(n58), .CP(clk), .CDN(rst_n), .Q(Q_mag[9]) );
  DFCNQD1 \Q_mag_reg[5]  ( .D(n62), .CP(clk), .CDN(rst_n), .Q(Q_mag[5]) );
  DFCNQD1 \Q_mag_reg[21]  ( .D(n46), .CP(clk), .CDN(rst_n), .Q(Q_mag[21]) );
  DFCNQD1 \Q_mag_reg[1]  ( .D(n66), .CP(clk), .CDN(rst_n), .Q(Q_mag[1]) );
  DFCNQD1 \Q_mag_reg[17]  ( .D(n50), .CP(clk), .CDN(rst_n), .Q(Q_mag[17]) );
  DFCNQD1 \Q_mag_reg[13]  ( .D(n54), .CP(clk), .CDN(rst_n), .Q(Q_mag[13]) );
  DFCNQD1 \Q_mag_reg[7]  ( .D(n60), .CP(clk), .CDN(rst_n), .Q(Q_mag[7]) );
  DFCNQD1 \Q_mag_reg[3]  ( .D(n64), .CP(clk), .CDN(rst_n), .Q(Q_mag[3]) );
  DFCNQD1 \Q_mag_reg[19]  ( .D(n48), .CP(clk), .CDN(rst_n), .Q(Q_mag[19]) );
  DFCNQD1 \Q_mag_reg[15]  ( .D(n52), .CP(clk), .CDN(rst_n), .Q(Q_mag[15]) );
  DFCNQD1 \Q_mag_reg[11]  ( .D(n56), .CP(clk), .CDN(rst_n), .Q(Q_mag[11]) );
  DFCNQD1 \Q_mag_reg[6]  ( .D(n61), .CP(clk), .CDN(rst_n), .Q(Q_mag[6]) );
  DFCNQD1 \Q_mag_reg[2]  ( .D(n65), .CP(clk), .CDN(rst_n), .Q(Q_mag[2]) );
  DFCNQD1 \Q_mag_reg[22]  ( .D(n68), .CP(clk), .CDN(rst_n), .Q(Q_mag[22]) );
  DFCNQD1 \Q_mag_reg[18]  ( .D(n49), .CP(clk), .CDN(rst_n), .Q(Q_mag[18]) );
  DFCNQD1 \Q_mag_reg[14]  ( .D(n53), .CP(clk), .CDN(rst_n), .Q(Q_mag[14]) );
  DFCNQD1 \Q_mag_reg[10]  ( .D(n57), .CP(clk), .CDN(rst_n), .Q(Q_mag[10]) );
  DFCNQD1 \Q_mag_reg[8]  ( .D(n59), .CP(clk), .CDN(rst_n), .Q(Q_mag[8]) );
  DFCNQD1 \Q_mag_reg[4]  ( .D(n63), .CP(clk), .CDN(rst_n), .Q(Q_mag[4]) );
  DFCNQD1 \Q_mag_reg[20]  ( .D(n47), .CP(clk), .CDN(rst_n), .Q(Q_mag[20]) );
  DFCNQD1 \Q_mag_reg[16]  ( .D(n51), .CP(clk), .CDN(rst_n), .Q(Q_mag[16]) );
  DFCNQD1 \Q_mag_reg[12]  ( .D(n55), .CP(clk), .CDN(rst_n), .Q(Q_mag[12]) );
  DFCNQD1 \Q_mag_reg[0]  ( .D(n67), .CP(clk), .CDN(rst_n), .Q(Q_mag[0]) );
  AO21D0 U3 ( .A1(n1017), .A2(n1027), .B(Q_mag[20]), .Z(n644) );
  INVD0 U4 ( .I(n644), .ZN(n600) );
  AO21D0 U5 ( .A1(n1019), .A2(n1017), .B(Q_mag[8]), .Z(n927) );
  INVD0 U6 ( .I(n927), .ZN(n839) );
  INVD0 U7 ( .I(n1030), .ZN(n828) );
  INVD0 U8 ( .I(n1029), .ZN(n698) );
  INVD0 U9 ( .I(n1028), .ZN(n1001) );
  AO21D0 U10 ( .A1(n1020), .A2(n1012), .B(Q_mag[14]), .Z(n774) );
  INVD0 U11 ( .I(n774), .ZN(n709) );
  AO21D0 U12 ( .A1(n1012), .A2(n1015), .B(Q_mag[2]), .Z(n1031) );
  INVD0 U13 ( .I(n1031), .ZN(n1032) );
  AOI22D0 U14 ( .A1(S_mag[3]), .A2(n702), .B1(S_mag[4]), .B2(n701), .ZN(n457)
         );
  NR2D0 U15 ( .A1(n902), .A2(n767), .ZN(n756) );
  NR2D0 U16 ( .A1(n882), .A2(n920), .ZN(n876) );
  NR2D0 U17 ( .A1(n919), .A2(n637), .ZN(n641) );
  NR2D0 U18 ( .A1(n919), .A2(n767), .ZN(n765) );
  AOI22D0 U19 ( .A1(S_mag[12]), .A2(n831), .B1(n977), .B2(n829), .ZN(n811) );
  OAI22D0 U20 ( .A1(n917), .A2(n638), .B1(n919), .B2(n639), .ZN(n634) );
  OAI22D0 U21 ( .A1(n911), .A2(n769), .B1(n902), .B2(n768), .ZN(n758) );
  NR2D0 U22 ( .A1(n911), .A2(n767), .ZN(n762) );
  AOI22D0 U23 ( .A1(n1006), .A2(S_mag[8]), .B1(n1005), .B2(S_mag[7]), .ZN(n994) );
  INVD0 U24 ( .I(n548), .ZN(\DP_OP_13J3_123_8774/n546 ) );
  AOI22D0 U25 ( .A1(S_mag[13]), .A2(n700), .B1(n965), .B2(n699), .ZN(n672) );
  AOI211D0 U26 ( .A1(n642), .A2(n981), .B(n494), .C(n493), .ZN(n495) );
  AOI22D0 U27 ( .A1(n179), .A2(S_mag[11]), .B1(n178), .B2(S_mag[10]), .ZN(n150) );
  NR2D0 U28 ( .A1(n886), .A2(n916), .ZN(n884) );
  CKND2D0 U29 ( .A1(n955), .A2(n954), .ZN(n956) );
  NR2D0 U30 ( .A1(n906), .A2(n916), .ZN(n904) );
  AOI211D0 U31 ( .A1(n772), .A2(n985), .B(n747), .C(n746), .ZN(n748) );
  OAI22D0 U32 ( .A1(n911), .A2(n638), .B1(n906), .B2(n639), .ZN(n628) );
  OAI22D0 U33 ( .A1(n930), .A2(n768), .B1(n769), .B2(n850), .ZN(n713) );
  AOI22D0 U34 ( .A1(S_mag[14]), .A2(n701), .B1(S_mag[13]), .B2(n702), .ZN(n674) );
  OAI22D0 U35 ( .A1(n870), .A2(n584), .B1(n866), .B2(n585), .ZN(n488) );
  AOI22D0 U36 ( .A1(n1006), .A2(S_mag[4]), .B1(n1005), .B2(S_mag[3]), .ZN(n90)
         );
  AOI22D0 U37 ( .A1(n177), .A2(S_mag[16]), .B1(n176), .B2(n953), .ZN(n21) );
  AOI22D0 U38 ( .A1(n1006), .A2(S_mag[20]), .B1(n1005), .B2(S_mag[19]), .ZN(
        n946) );
  AOI21D0 U39 ( .A1(n1020), .A2(n446), .B(Q_mag[15]), .ZN(n451) );
  AOI211D0 U40 ( .A1(n981), .A2(n772), .B(n744), .C(n743), .ZN(n745) );
  CKND2D0 U41 ( .A1(n544), .A2(n543), .ZN(\DP_OP_13J3_123_8774/n737 ) );
  AOI21D0 U42 ( .A1(n1019), .A2(n1013), .B(Q_mag[9]), .ZN(n420) );
  OAI22D0 U43 ( .A1(n933), .A2(n778), .B1(n928), .B2(n776), .ZN(n775) );
  AOI211D0 U44 ( .A1(n772), .A2(n937), .B(n711), .C(n710), .ZN(n712) );
  AOI22D0 U45 ( .A1(S_mag[11]), .A2(n571), .B1(n570), .B2(n981), .ZN(n533) );
  CKND2D0 U46 ( .A1(n113), .A2(n112), .ZN(n114) );
  AOI22D0 U47 ( .A1(n179), .A2(S_mag[12]), .B1(n176), .B2(n977), .ZN(n37) );
  CKND2D0 U48 ( .A1(n947), .A2(n946), .ZN(n948) );
  AOI22D0 U49 ( .A1(n178), .A2(S_mag[12]), .B1(n177), .B2(S_mag[11]), .ZN(n155) );
  INVD0 U50 ( .I(S_mag[1]), .ZN(n921) );
  AOI21D0 U51 ( .A1(n1018), .A2(n1017), .B(Q_mag[4]), .ZN(n76) );
  CKND2D0 U52 ( .A1(n526), .A2(n525), .ZN(\DP_OP_13J3_123_8774/n736 ) );
  INVD0 U53 ( .I(n646), .ZN(n699) );
  INVD0 U54 ( .I(\DP_OP_13J3_123_8774/n436 ), .ZN(n358) );
  INVD0 U55 ( .I(n498), .ZN(\DP_OP_13J3_123_8774/n466 ) );
  AOI22D0 U56 ( .A1(n179), .A2(S_mag[7]), .B1(n178), .B2(S_mag[6]), .ZN(n131)
         );
  INVD0 U57 ( .I(n205), .ZN(n206) );
  AOI211D0 U58 ( .A1(n925), .A2(n993), .B(n896), .C(n895), .ZN(n897) );
  CKND2D0 U59 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  AOI211D0 U60 ( .A1(n642), .A2(n985), .B(n617), .C(n616), .ZN(n618) );
  CKND2D0 U61 ( .A1(n939), .A2(n938), .ZN(n940) );
  CKND2D0 U62 ( .A1(n684), .A2(n683), .ZN(n685) );
  INVD0 U63 ( .I(\DP_OP_13J3_123_8774/n435 ), .ZN(n349) );
  CKND2D0 U64 ( .A1(n370), .A2(n367), .ZN(n365) );
  CKND2D0 U65 ( .A1(n528), .A2(n527), .ZN(\DP_OP_13J3_123_8774/n723 ) );
  CKND2D0 U66 ( .A1(n127), .A2(n126), .ZN(n128) );
  OAI22D0 U67 ( .A1(n211), .A2(n210), .B1(n208), .B2(n209), .ZN(n207) );
  AOI22D0 U68 ( .A1(n179), .A2(S_mag[15]), .B1(n178), .B2(S_mag[14]), .ZN(n28)
         );
  CKND2D0 U69 ( .A1(n33), .A2(n32), .ZN(n34) );
  INVD0 U70 ( .I(n299), .ZN(n142) );
  CKND2D0 U71 ( .A1(n83), .A2(n78), .ZN(n934) );
  CKND2D0 U72 ( .A1(n514), .A2(n513), .ZN(\DP_OP_13J3_123_8774/n733 ) );
  INVD0 U73 ( .I(n348), .ZN(n355) );
  NR2D0 U74 ( .A1(n311), .A2(n310), .ZN(n573) );
  AOI22D0 U75 ( .A1(S_mag[20]), .A2(n573), .B1(n937), .B2(n570), .ZN(n312) );
  CKND2D0 U76 ( .A1(n281), .A2(n280), .ZN(n288) );
  AOI211D0 U77 ( .A1(n925), .A2(n937), .B(n841), .C(n840), .ZN(n842) );
  CKND2D0 U78 ( .A1(n793), .A2(n792), .ZN(n794) );
  OAI21D0 U79 ( .A1(n381), .A2(n380), .B(n379), .ZN(n386) );
  OAI21D0 U80 ( .A1(n600), .A2(\DP_OP_13J3_123_8774/n388 ), .B(n327), .ZN(n388) );
  AOI32D0 U81 ( .A1(n388), .A2(n335), .A3(n389), .B1(n387), .B2(n335), .ZN(
        n396) );
  CKND2D0 U82 ( .A1(n402), .A2(n401), .ZN(n562) );
  OAI21D0 U83 ( .A1(n403), .A2(n406), .B(n562), .ZN(n69) );
  NR2D0 U84 ( .A1(bit_pos[1]), .A2(bit_pos[0]), .ZN(n1017) );
  INVD0 U85 ( .I(bit_pos[2]), .ZN(n407) );
  CKND2D0 U86 ( .A1(n1017), .A2(n407), .ZN(n1) );
  NR2D0 U87 ( .A1(bit_pos[3]), .A2(n1), .ZN(n402) );
  INVD0 U88 ( .I(bit_pos[4]), .ZN(n305) );
  CKND2D0 U89 ( .A1(n402), .A2(n305), .ZN(n405) );
  CKND2D0 U90 ( .A1(running), .A2(n405), .ZN(n1011) );
  INVD0 U91 ( .I(n1011), .ZN(n401) );
  CKND2D0 U92 ( .A1(n1017), .A2(n401), .ZN(n2) );
  INVD0 U93 ( .I(running), .ZN(n404) );
  CKND2D0 U94 ( .A1(start), .A2(n404), .ZN(n1025) );
  OAI21D0 U95 ( .A1(n1), .A2(n1011), .B(n1025), .ZN(n403) );
  AO21D0 U96 ( .A1(bit_pos[2]), .A2(n2), .B(n403), .Z(n70) );
  INVD0 U97 ( .I(n1025), .ZN(n400) );
  AOI221D0 U98 ( .A1(n1017), .A2(n401), .B1(bit_pos[1]), .B2(n1011), .C(n400), 
        .ZN(n3) );
  CKND2D0 U99 ( .A1(bit_pos[1]), .A2(bit_pos[0]), .ZN(n1014) );
  CKND2D0 U100 ( .A1(n3), .A2(n1014), .ZN(n71) );
  INVD0 U101 ( .I(bit_pos[0]), .ZN(n1010) );
  NR2D0 U102 ( .A1(bit_pos[1]), .A2(n1010), .ZN(n1013) );
  INVD0 U103 ( .I(bit_pos[3]), .ZN(n406) );
  CKND2D0 U104 ( .A1(bit_pos[2]), .A2(n406), .ZN(n306) );
  NR2D0 U105 ( .A1(bit_pos[4]), .A2(n306), .ZN(n1018) );
  AOI21D1 U106 ( .A1(n1013), .A2(n1018), .B(Q_mag[5]), .ZN(n1028) );
  NR3D0 U107 ( .A1(bit_pos[2]), .A2(bit_pos[4]), .A3(n406), .ZN(n1019) );
  INVD0 U108 ( .I(n1014), .ZN(n446) );
  AOI21D1 U109 ( .A1(n1019), .A2(n446), .B(Q_mag[11]), .ZN(n1030) );
  INR2D0 U110 ( .A1(bit_pos[1]), .B1(bit_pos[0]), .ZN(n1012) );
  NR3D0 U111 ( .A1(bit_pos[3]), .A2(bit_pos[2]), .A3(bit_pos[4]), .ZN(n1015)
         );
  NR3D0 U112 ( .A1(bit_pos[3]), .A2(bit_pos[2]), .A3(n305), .ZN(n1023) );
  AOI21D1 U113 ( .A1(n1023), .A2(n1013), .B(Q_mag[17]), .ZN(n1029) );
  AOI21D0 U114 ( .A1(n446), .A2(n1018), .B(Q_mag[7]), .ZN(n4) );
  MUX2ND0 U115 ( .I0(n927), .I1(n839), .S(n4), .ZN(n9) );
  AOI21D0 U116 ( .A1(n1018), .A2(n1012), .B(Q_mag[6]), .ZN(n6) );
  INVD0 U117 ( .I(n6), .ZN(n5) );
  MUX2ND0 U118 ( .I0(n1028), .I1(n1001), .S(n5), .ZN(n10) );
  IND2D0 U119 ( .A1(n9), .B1(n10), .ZN(n918) );
  INVD0 U120 ( .I(S_mag[0]), .ZN(n583) );
  MUX2ND0 U121 ( .I0(n6), .I1(n5), .S(n4), .ZN(n8) );
  OR2D0 U122 ( .A1(n8), .A2(n10), .Z(n916) );
  OAI22D0 U123 ( .A1(n921), .A2(S_mag[0]), .B1(n583), .B2(S_mag[1]), .ZN(n462)
         );
  INVD0 U124 ( .I(n462), .ZN(n586) );
  CKND2D0 U125 ( .A1(n10), .A2(n9), .ZN(n837) );
  OA222D0 U126 ( .A1(n921), .A2(n918), .B1(n583), .B2(n916), .C1(n586), .C2(
        n837), .Z(n94) );
  CKND2D0 U127 ( .A1(S_mag[0]), .A2(n10), .ZN(n122) );
  ND3D0 U128 ( .A1(n94), .A2(n122), .A3(n927), .ZN(n44) );
  INVD0 U129 ( .I(n837), .ZN(n925) );
  INVD0 U130 ( .I(S_mag[2]), .ZN(n917) );
  NR2D0 U131 ( .A1(S_mag[0]), .A2(n921), .ZN(n7) );
  MUX2ND0 U132 ( .I0(n917), .I1(S_mag[2]), .S(n7), .ZN(n542) );
  NR2D0 U133 ( .A1(n921), .A2(n916), .ZN(n12) );
  IND3D0 U134 ( .A1(n10), .B1(n9), .B2(n8), .ZN(n920) );
  OAI22D0 U135 ( .A1(n917), .A2(n918), .B1(n583), .B2(n920), .ZN(n11) );
  AOI211D0 U136 ( .A1(n925), .A2(n542), .B(n12), .C(n11), .ZN(n45) );
  CKND2D0 U137 ( .A1(n45), .A2(n927), .ZN(n43) );
  NR2D0 U138 ( .A1(n44), .A2(n43), .ZN(\DP_OP_13J3_123_8774/n631 ) );
  INVD0 U139 ( .I(Q_mag[0]), .ZN(n399) );
  AOI21D0 U140 ( .A1(n917), .A2(n583), .B(n921), .ZN(n85) );
  CKND2D0 U141 ( .A1(S_mag[22]), .A2(n13), .ZN(n928) );
  OAI21D0 U142 ( .A1(S_mag[22]), .A2(n13), .B(n928), .ZN(n935) );
  CKND2D0 U143 ( .A1(n399), .A2(n405), .ZN(n18) );
  AOI21D0 U144 ( .A1(n1015), .A2(n1013), .B(Q_mag[1]), .ZN(n14) );
  MUX2ND0 U145 ( .I0(n1031), .I1(n1032), .S(n14), .ZN(n19) );
  CKND2D0 U146 ( .A1(n18), .A2(n19), .ZN(n184) );
  INVD0 U147 ( .I(S_mag[22]), .ZN(n933) );
  NR2D0 U148 ( .A1(n14), .A2(n18), .ZN(n178) );
  INVD0 U149 ( .I(n178), .ZN(n104) );
  CKND2D0 U150 ( .A1(n14), .A2(n1031), .ZN(n15) );
  NR2D0 U151 ( .A1(n18), .A2(n15), .ZN(n177) );
  INVD0 U152 ( .I(n177), .ZN(n185) );
  INVD0 U153 ( .I(S_mag[21]), .ZN(n930) );
  OAI222D0 U154 ( .A1(n935), .A2(n184), .B1(n933), .B2(n104), .C1(n185), .C2(
        n930), .ZN(n16) );
  MUX2ND0 U155 ( .I0(n1032), .I1(n1031), .S(n16), .ZN(n202) );
  INVD0 U156 ( .I(\DP_OP_13J3_123_8774/n532 ), .ZN(n225) );
  INVD0 U157 ( .I(\DP_OP_13J3_123_8774/n541 ), .ZN(n222) );
  INVD0 U158 ( .I(\DP_OP_13J3_123_8774/n551 ), .ZN(n235) );
  INVD0 U159 ( .I(n184), .ZN(n176) );
  FA1D0 U160 ( .A(S_mag[17]), .B(S_mag[18]), .CI(n17), .CO(n163), .S(n953) );
  INVD0 U161 ( .I(n18), .ZN(n105) );
  NR2D0 U162 ( .A1(n105), .A2(n19), .ZN(n179) );
  AOI22D0 U163 ( .A1(n179), .A2(S_mag[18]), .B1(n178), .B2(S_mag[17]), .ZN(n20) );
  CKND2D0 U164 ( .A1(n21), .A2(n20), .ZN(n22) );
  MUX2ND0 U165 ( .I0(n1032), .I1(n1031), .S(n22), .ZN(n196) );
  FA1D0 U166 ( .A(S_mag[16]), .B(S_mag[17]), .CI(n23), .CO(n17), .S(n957) );
  AOI22D0 U167 ( .A1(n177), .A2(S_mag[15]), .B1(n176), .B2(n957), .ZN(n25) );
  AOI22D0 U168 ( .A1(n179), .A2(S_mag[17]), .B1(n178), .B2(S_mag[16]), .ZN(n24) );
  CKND2D0 U169 ( .A1(n25), .A2(n24), .ZN(n26) );
  MUX2ND0 U170 ( .I0(n1032), .I1(n1031), .S(n26), .ZN(n209) );
  INVD0 U171 ( .I(\DP_OP_13J3_123_8774/n579 ), .ZN(n228) );
  FA1D0 U172 ( .A(S_mag[14]), .B(S_mag[15]), .CI(n27), .CO(n158), .S(n965) );
  AOI22D0 U173 ( .A1(n177), .A2(S_mag[13]), .B1(n176), .B2(n965), .ZN(n29) );
  CKND2D0 U174 ( .A1(n29), .A2(n28), .ZN(n30) );
  MUX2ND0 U175 ( .I0(n1032), .I1(n1031), .S(n30), .ZN(n190) );
  FA1D0 U176 ( .A(S_mag[13]), .B(S_mag[14]), .CI(n31), .CO(n27), .S(n969) );
  AOI22D0 U177 ( .A1(n177), .A2(S_mag[12]), .B1(n176), .B2(n969), .ZN(n33) );
  AOI22D0 U178 ( .A1(n179), .A2(S_mag[14]), .B1(n178), .B2(S_mag[13]), .ZN(n32) );
  MUX2ND0 U179 ( .I0(n1031), .I1(n1032), .S(n34), .ZN(n277) );
  INVD0 U180 ( .I(\DP_OP_13J3_123_8774/n595 ), .ZN(n274) );
  FA1D0 U181 ( .A(S_mag[11]), .B(S_mag[12]), .CI(n35), .CO(n154), .S(n977) );
  AOI22D0 U182 ( .A1(n178), .A2(S_mag[11]), .B1(n177), .B2(S_mag[10]), .ZN(n36) );
  CKND2D0 U183 ( .A1(n37), .A2(n36), .ZN(n38) );
  MUX2ND0 U184 ( .I0(n1032), .I1(n1031), .S(n38), .ZN(n211) );
  INVD0 U185 ( .I(\DP_OP_13J3_123_8774/n616 ), .ZN(n238) );
  FA1D0 U186 ( .A(S_mag[9]), .B(S_mag[10]), .CI(n39), .CO(n149), .S(n985) );
  AOI22D0 U187 ( .A1(n177), .A2(S_mag[8]), .B1(n176), .B2(n985), .ZN(n41) );
  AOI22D0 U188 ( .A1(n179), .A2(S_mag[10]), .B1(n178), .B2(S_mag[9]), .ZN(n40)
         );
  CKND2D0 U189 ( .A1(n41), .A2(n40), .ZN(n42) );
  MUX2ND0 U190 ( .I0(n1032), .I1(n1031), .S(n42), .ZN(n188) );
  OAI211D0 U191 ( .A1(n45), .A2(n927), .B(n44), .C(n43), .ZN(n75) );
  IND2D0 U192 ( .A1(\DP_OP_13J3_123_8774/n631 ), .B1(n75), .ZN(n475) );
  MUX2ND0 U193 ( .I0(n1001), .I1(n1028), .S(n76), .ZN(n78) );
  AOI21D0 U194 ( .A1(n1015), .A2(n446), .B(Q_mag[3]), .ZN(n77) );
  CKXOR2D0 U195 ( .A1(n77), .A2(n76), .Z(n80) );
  MUX2ND0 U196 ( .I0(n1031), .I1(n1032), .S(n77), .ZN(n83) );
  INR3D0 U197 ( .A1(n78), .B1(n80), .B2(n83), .ZN(n1004) );
  INVD0 U198 ( .I(n934), .ZN(n1003) );
  AOI22D0 U199 ( .A1(S_mag[0]), .A2(n1004), .B1(n1003), .B2(n542), .ZN(n82) );
  INVD0 U200 ( .I(n83), .ZN(n79) );
  NR2D0 U201 ( .A1(n79), .A2(n78), .ZN(n1006) );
  CKND2D0 U202 ( .A1(n80), .A2(n79), .ZN(n932) );
  INVD0 U203 ( .I(n932), .ZN(n1005) );
  AOI22D0 U204 ( .A1(n1006), .A2(S_mag[2]), .B1(S_mag[1]), .B2(n1005), .ZN(n81) );
  CKND2D0 U205 ( .A1(n82), .A2(n81), .ZN(n101) );
  INVD0 U206 ( .I(n101), .ZN(n84) );
  CKND2D0 U207 ( .A1(n83), .A2(S_mag[0]), .ZN(n111) );
  AOI222D0 U208 ( .A1(S_mag[0]), .A2(n1005), .B1(S_mag[1]), .B2(n1006), .C1(
        n1003), .C2(n462), .ZN(n103) );
  AN3D0 U209 ( .A1(n1001), .A2(n111), .A3(n103), .Z(n100) );
  CKND2D0 U210 ( .A1(n84), .A2(n100), .ZN(n123) );
  FA1D0 U211 ( .A(S_mag[2]), .B(S_mag[3]), .CI(n85), .CO(n89), .S(n924) );
  AOI22D0 U212 ( .A1(S_mag[1]), .A2(n1004), .B1(n1003), .B2(n924), .ZN(n87) );
  AOI22D0 U213 ( .A1(n1006), .A2(S_mag[3]), .B1(S_mag[2]), .B2(n1005), .ZN(n86) );
  CKND2D0 U214 ( .A1(n87), .A2(n86), .ZN(n88) );
  MUX2ND0 U215 ( .I0(n1028), .I1(n1001), .S(n88), .ZN(n124) );
  IOA21D0 U216 ( .A1(n123), .A2(n122), .B(n124), .ZN(n136) );
  FA1D0 U217 ( .A(S_mag[3]), .B(S_mag[4]), .CI(n89), .CO(n95), .S(n914) );
  AOI22D0 U218 ( .A1(S_mag[2]), .A2(n1004), .B1(n1003), .B2(n914), .ZN(n91) );
  CKND2D0 U219 ( .A1(n91), .A2(n90), .ZN(n92) );
  MUX2ND0 U220 ( .I0(n1001), .I1(n1028), .S(n92), .ZN(n135) );
  OAI21D0 U221 ( .A1(n839), .A2(n122), .B(n94), .ZN(n93) );
  OAI31D0 U222 ( .A1(n839), .A2(n94), .A3(n122), .B(n93), .ZN(n134) );
  FA1D0 U223 ( .A(S_mag[4]), .B(S_mag[5]), .CI(n95), .CO(n125), .S(n909) );
  AOI22D0 U224 ( .A1(n1004), .A2(S_mag[3]), .B1(n1003), .B2(n909), .ZN(n97) );
  AOI22D0 U225 ( .A1(n1006), .A2(S_mag[5]), .B1(n1005), .B2(S_mag[4]), .ZN(n96) );
  CKND2D0 U226 ( .A1(n97), .A2(n96), .ZN(n98) );
  MUX2ND0 U227 ( .I0(n1001), .I1(n1028), .S(n98), .ZN(n473) );
  MAOI222D0 U228 ( .A(n101), .B(n100), .C(n1028), .ZN(n99) );
  OAI31D0 U229 ( .A1(n101), .A2(n100), .A3(n1028), .B(n99), .ZN(n272) );
  OAI21D0 U230 ( .A1(n1028), .A2(n111), .B(n103), .ZN(n102) );
  OA31D0 U231 ( .A1(n1028), .A2(n103), .A3(n111), .B(n102), .Z(n258) );
  OAI222D0 U232 ( .A1(n105), .A2(n921), .B1(n105), .B2(n583), .C1(n583), .C2(
        n104), .ZN(n214) );
  NR2D0 U233 ( .A1(n1032), .A2(n214), .ZN(n109) );
  AOI22D0 U234 ( .A1(S_mag[0]), .A2(n177), .B1(n542), .B2(n176), .ZN(n107) );
  AOI22D0 U235 ( .A1(S_mag[2]), .A2(n179), .B1(S_mag[1]), .B2(n178), .ZN(n106)
         );
  CKND2D0 U236 ( .A1(n107), .A2(n106), .ZN(n257) );
  INVD0 U237 ( .I(n257), .ZN(n108) );
  CKND2D0 U238 ( .A1(n109), .A2(n108), .ZN(n110) );
  CKND2D0 U239 ( .A1(n111), .A2(n110), .ZN(n255) );
  AOI22D0 U240 ( .A1(S_mag[1]), .A2(n177), .B1(n176), .B2(n924), .ZN(n113) );
  AOI22D0 U241 ( .A1(S_mag[2]), .A2(n178), .B1(n179), .B2(S_mag[3]), .ZN(n112)
         );
  MUX2ND0 U242 ( .I0(n1031), .I1(n1032), .S(n114), .ZN(n254) );
  INR2D0 U243 ( .A1(n255), .B1(n254), .ZN(n259) );
  AOI22D0 U244 ( .A1(S_mag[2]), .A2(n177), .B1(n176), .B2(n914), .ZN(n116) );
  AOI22D0 U245 ( .A1(n179), .A2(S_mag[4]), .B1(S_mag[3]), .B2(n178), .ZN(n115)
         );
  CKND2D0 U246 ( .A1(n116), .A2(n115), .ZN(n117) );
  MUX2ND0 U247 ( .I0(n1032), .I1(n1031), .S(n117), .ZN(n265) );
  MAOI222D0 U248 ( .A(n258), .B(n259), .C(n265), .ZN(n118) );
  INVD0 U249 ( .I(n118), .ZN(n271) );
  AOI22D0 U250 ( .A1(S_mag[3]), .A2(n177), .B1(n176), .B2(n909), .ZN(n120) );
  AOI22D0 U251 ( .A1(n179), .A2(S_mag[5]), .B1(n178), .B2(S_mag[4]), .ZN(n119)
         );
  CKND2D0 U252 ( .A1(n120), .A2(n119), .ZN(n121) );
  MUX2ND0 U253 ( .I0(n1032), .I1(n1031), .S(n121), .ZN(n278) );
  MAOI222D0 U254 ( .A(n272), .B(n271), .C(n278), .ZN(n283) );
  XNR3D0 U255 ( .A1(n124), .A2(n123), .A3(n122), .ZN(n282) );
  FA1D0 U256 ( .A(S_mag[5]), .B(S_mag[6]), .CI(n125), .CO(n130), .S(n1002) );
  AOI22D0 U257 ( .A1(n177), .A2(S_mag[4]), .B1(n176), .B2(n1002), .ZN(n127) );
  AOI22D0 U258 ( .A1(n179), .A2(S_mag[6]), .B1(n178), .B2(S_mag[5]), .ZN(n126)
         );
  MUX2ND0 U259 ( .I0(n1031), .I1(n1032), .S(n128), .ZN(n285) );
  MAOI222D0 U260 ( .A(n283), .B(n282), .C(n285), .ZN(n129) );
  INVD0 U261 ( .I(n129), .ZN(n280) );
  FA1D0 U262 ( .A(S_mag[6]), .B(S_mag[7]), .CI(n130), .CO(n138), .S(n997) );
  AOI22D0 U263 ( .A1(n177), .A2(S_mag[5]), .B1(n176), .B2(n997), .ZN(n132) );
  CKND2D0 U264 ( .A1(n132), .A2(n131), .ZN(n133) );
  MUX2ND0 U265 ( .I0(n1031), .I1(n1032), .S(n133), .ZN(n287) );
  FA1D0 U266 ( .A(n136), .B(n135), .CI(n134), .CO(n474), .S(n281) );
  MAOI222D0 U267 ( .A(n280), .B(n287), .C(n281), .ZN(n137) );
  INVD0 U268 ( .I(n137), .ZN(n295) );
  FA1D0 U269 ( .A(S_mag[7]), .B(S_mag[8]), .CI(n138), .CO(n143), .S(n993) );
  AOI22D0 U270 ( .A1(n177), .A2(S_mag[6]), .B1(n176), .B2(n993), .ZN(n140) );
  AOI22D0 U271 ( .A1(n179), .A2(S_mag[8]), .B1(n178), .B2(S_mag[7]), .ZN(n139)
         );
  CKND2D0 U272 ( .A1(n140), .A2(n139), .ZN(n141) );
  MUX2ND0 U273 ( .I0(n1032), .I1(n1031), .S(n141), .ZN(n299) );
  MAOI222D0 U274 ( .A(n296), .B(n295), .C(n142), .ZN(n147) );
  FA1D0 U275 ( .A(S_mag[8]), .B(S_mag[9]), .CI(n143), .CO(n39), .S(n989) );
  AOI22D0 U276 ( .A1(n177), .A2(S_mag[7]), .B1(n176), .B2(n989), .ZN(n145) );
  AOI22D0 U277 ( .A1(n179), .A2(S_mag[9]), .B1(n178), .B2(S_mag[8]), .ZN(n144)
         );
  CKND2D0 U278 ( .A1(n145), .A2(n144), .ZN(n146) );
  MUX2ND0 U279 ( .I0(n1032), .I1(n1031), .S(n146), .ZN(n293) );
  MAOI222D0 U280 ( .A(n147), .B(n293), .C(\DP_OP_13J3_123_8774/n626 ), .ZN(
        n189) );
  INVD0 U281 ( .I(n189), .ZN(n148) );
  MAOI222D0 U282 ( .A(\DP_OP_13J3_123_8774/n621 ), .B(n188), .C(n148), .ZN(
        n237) );
  FA1D0 U283 ( .A(S_mag[10]), .B(S_mag[11]), .CI(n149), .CO(n35), .S(n981) );
  AOI22D0 U284 ( .A1(n177), .A2(S_mag[9]), .B1(n176), .B2(n981), .ZN(n151) );
  CKND2D0 U285 ( .A1(n151), .A2(n150), .ZN(n152) );
  MUX2ND0 U286 ( .I0(n1031), .I1(n1032), .S(n152), .ZN(n236) );
  INVD0 U287 ( .I(n203), .ZN(n204) );
  MAOI222D0 U288 ( .A(n211), .B(\DP_OP_13J3_123_8774/n609 ), .C(n204), .ZN(
        n153) );
  INVD0 U289 ( .I(n153), .ZN(n260) );
  FA1D0 U290 ( .A(S_mag[12]), .B(S_mag[13]), .CI(n154), .CO(n31), .S(n973) );
  AOI22D0 U291 ( .A1(n179), .A2(S_mag[13]), .B1(n176), .B2(n973), .ZN(n156) );
  CKND2D0 U292 ( .A1(n156), .A2(n155), .ZN(n157) );
  MUX2ND0 U293 ( .I0(n1032), .I1(n1031), .S(n157), .ZN(n263) );
  MAOI222D0 U294 ( .A(n260), .B(n263), .C(\DP_OP_13J3_123_8774/n602 ), .ZN(
        n273) );
  MAOI222D0 U295 ( .A(n277), .B(n274), .C(n273), .ZN(n191) );
  MAOI222D0 U296 ( .A(\DP_OP_13J3_123_8774/n587 ), .B(n190), .C(n191), .ZN(
        n227) );
  FA1D0 U297 ( .A(S_mag[15]), .B(S_mag[16]), .CI(n158), .CO(n23), .S(n961) );
  AOI22D0 U298 ( .A1(n177), .A2(S_mag[14]), .B1(n176), .B2(n961), .ZN(n160) );
  AOI22D0 U299 ( .A1(n179), .A2(S_mag[16]), .B1(n178), .B2(S_mag[15]), .ZN(
        n159) );
  CKND2D0 U300 ( .A1(n160), .A2(n159), .ZN(n161) );
  MUX2ND0 U301 ( .I0(n1031), .I1(n1032), .S(n161), .ZN(n226) );
  MAOI222D0 U302 ( .A(n209), .B(\DP_OP_13J3_123_8774/n571 ), .C(n206), .ZN(
        n200) );
  INVD0 U303 ( .I(n200), .ZN(n162) );
  MAOI222D0 U304 ( .A(\DP_OP_13J3_123_8774/n561 ), .B(n196), .C(n162), .ZN(
        n234) );
  FA1D0 U305 ( .A(S_mag[18]), .B(S_mag[19]), .CI(n163), .CO(n167), .S(n949) );
  AOI22D0 U306 ( .A1(n177), .A2(S_mag[17]), .B1(n176), .B2(n949), .ZN(n165) );
  AOI22D0 U307 ( .A1(n179), .A2(S_mag[19]), .B1(n178), .B2(S_mag[18]), .ZN(
        n164) );
  CKND2D0 U308 ( .A1(n165), .A2(n164), .ZN(n166) );
  MUX2ND0 U309 ( .I0(n1031), .I1(n1032), .S(n166), .ZN(n233) );
  FA1D0 U310 ( .A(S_mag[19]), .B(S_mag[20]), .CI(n167), .CO(n171), .S(n945) );
  AOI22D0 U311 ( .A1(n177), .A2(S_mag[18]), .B1(n176), .B2(n945), .ZN(n169) );
  AOI22D0 U312 ( .A1(n179), .A2(S_mag[20]), .B1(n178), .B2(S_mag[19]), .ZN(
        n168) );
  CKND2D0 U313 ( .A1(n169), .A2(n168), .ZN(n170) );
  MUX2ND0 U314 ( .I0(n1031), .I1(n1032), .S(n170), .ZN(n220) );
  FA1D0 U315 ( .A(S_mag[20]), .B(S_mag[21]), .CI(n171), .CO(n175), .S(n941) );
  AOI22D0 U316 ( .A1(n177), .A2(S_mag[19]), .B1(n176), .B2(n941), .ZN(n173) );
  AOI22D0 U317 ( .A1(n179), .A2(S_mag[21]), .B1(n178), .B2(S_mag[20]), .ZN(
        n172) );
  CKND2D0 U318 ( .A1(n173), .A2(n172), .ZN(n174) );
  MUX2ND0 U319 ( .I0(n1031), .I1(n1032), .S(n174), .ZN(n223) );
  INVD0 U320 ( .I(n212), .ZN(n213) );
  FA1D0 U321 ( .A(S_mag[21]), .B(S_mag[22]), .CI(n175), .CO(n13), .S(n937) );
  AOI22D0 U322 ( .A1(n177), .A2(S_mag[20]), .B1(n176), .B2(n937), .ZN(n181) );
  AOI22D0 U323 ( .A1(n179), .A2(S_mag[22]), .B1(n178), .B2(S_mag[21]), .ZN(
        n180) );
  CKND2D0 U324 ( .A1(n181), .A2(n180), .ZN(n182) );
  MUX2ND0 U325 ( .I0(n1032), .I1(n1031), .S(n182), .ZN(n217) );
  MAOI222D0 U326 ( .A(n213), .B(n217), .C(\DP_OP_13J3_123_8774/n523 ), .ZN(
        n183) );
  INVD0 U327 ( .I(n183), .ZN(n194) );
  MAOI222D0 U328 ( .A(n202), .B(\DP_OP_13J3_123_8774/n514 ), .C(n194), .ZN(
        n193) );
  INVD0 U329 ( .I(\DP_OP_13J3_123_8774/n505 ), .ZN(n187) );
  OAI22D0 U330 ( .A1(n185), .A2(n933), .B1(n184), .B2(n928), .ZN(n186) );
  MUX2ND0 U331 ( .I0(n1031), .I1(n1032), .S(n186), .ZN(n192) );
  MAOI222D0 U332 ( .A(n193), .B(n187), .C(n192), .ZN(n219) );
  MAOI222D0 U333 ( .A(\DP_OP_13J3_123_8774/n487 ), .B(n240), .C(
        \DP_OP_13J3_123_8774/n495 ), .ZN(n244) );
  INVD0 U334 ( .I(\DP_OP_13J3_123_8774/n478 ), .ZN(n241) );
  INVD0 U335 ( .I(\DP_OP_13J3_123_8774/n486 ), .ZN(n242) );
  MAOI222D0 U336 ( .A(n244), .B(n241), .C(n242), .ZN(n324) );
  XOR3D0 U337 ( .A1(n189), .A2(\DP_OP_13J3_123_8774/n621 ), .A3(n188), .Z(n304) );
  XNR3D0 U338 ( .A1(n191), .A2(\DP_OP_13J3_123_8774/n587 ), .A3(n190), .ZN(
        n303) );
  XOR3D0 U339 ( .A1(n193), .A2(\DP_OP_13J3_123_8774/n505 ), .A3(n192), .Z(n292) );
  INVD0 U340 ( .I(\DP_OP_13J3_123_8774/n514 ), .ZN(n195) );
  MUX2ND0 U341 ( .I0(\DP_OP_13J3_123_8774/n514 ), .I1(n195), .S(n194), .ZN(
        n201) );
  INVD0 U342 ( .I(\DP_OP_13J3_123_8774/n561 ), .ZN(n197) );
  MUX2ND0 U343 ( .I0(n197), .I1(\DP_OP_13J3_123_8774/n561 ), .S(n196), .ZN(
        n199) );
  OAI22D0 U344 ( .A1(n202), .A2(n201), .B1(n199), .B2(n200), .ZN(n198) );
  AOI221D0 U345 ( .A1(n202), .A2(n201), .B1(n200), .B2(n199), .C(n198), .ZN(
        n270) );
  MUX2ND0 U346 ( .I0(n204), .I1(n203), .S(\DP_OP_13J3_123_8774/n609 ), .ZN(
        n210) );
  MUX2ND0 U347 ( .I0(n206), .I1(n205), .S(\DP_OP_13J3_123_8774/n571 ), .ZN(
        n208) );
  AOI221D0 U348 ( .A1(n211), .A2(n210), .B1(n209), .B2(n208), .C(n207), .ZN(
        n269) );
  MUX2ND0 U349 ( .I0(n213), .I1(n212), .S(\DP_OP_13J3_123_8774/n523 ), .ZN(
        n218) );
  INVD0 U350 ( .I(n214), .ZN(n215) );
  OAI21D0 U351 ( .A1(n218), .A2(n217), .B(n215), .ZN(n216) );
  AOI21D0 U352 ( .A1(n218), .A2(n217), .B(n216), .ZN(n253) );
  FA1D0 U353 ( .A(\DP_OP_13J3_123_8774/n504 ), .B(\DP_OP_13J3_123_8774/n496 ), 
        .CI(n219), .CO(n240), .S(n232) );
  FA1D0 U354 ( .A(n222), .B(n221), .CI(n220), .CO(n224), .S(n231) );
  FA1D0 U355 ( .A(n225), .B(n224), .CI(n223), .CO(n212), .S(n230) );
  FA1D0 U356 ( .A(n228), .B(n227), .CI(n226), .CO(n205), .S(n229) );
  IND4D0 U357 ( .A1(n232), .B1(n231), .B2(n230), .B3(n229), .ZN(n250) );
  FA1D0 U358 ( .A(n235), .B(n234), .CI(n233), .CO(n221), .S(n249) );
  FA1D0 U359 ( .A(n238), .B(n237), .CI(n236), .CO(n203), .S(n248) );
  INVD0 U360 ( .I(n240), .ZN(n239) );
  MUX2ND0 U361 ( .I0(n240), .I1(n239), .S(\DP_OP_13J3_123_8774/n495 ), .ZN(
        n246) );
  MUX2ND0 U362 ( .I0(\DP_OP_13J3_123_8774/n486 ), .I1(n242), .S(n241), .ZN(
        n245) );
  OAI22D0 U363 ( .A1(\DP_OP_13J3_123_8774/n487 ), .A2(n246), .B1(n245), .B2(
        n244), .ZN(n243) );
  AOI221D0 U364 ( .A1(n246), .A2(\DP_OP_13J3_123_8774/n487 ), .B1(n245), .B2(
        n244), .C(n243), .ZN(n247) );
  IND4D0 U365 ( .A1(n250), .B1(n249), .B2(n248), .B3(n247), .ZN(n251) );
  AOI21D0 U366 ( .A1(n255), .A2(n254), .B(n251), .ZN(n252) );
  OAI211D0 U367 ( .A1(n255), .A2(n254), .B(n253), .C(n252), .ZN(n256) );
  NR2D0 U368 ( .A1(n257), .A2(n256), .ZN(n268) );
  NR2D0 U369 ( .A1(n259), .A2(n258), .ZN(n266) );
  INVD0 U370 ( .I(\DP_OP_13J3_123_8774/n602 ), .ZN(n261) );
  MUX2ND0 U371 ( .I0(\DP_OP_13J3_123_8774/n602 ), .I1(n261), .S(n260), .ZN(
        n264) );
  OAI22D0 U372 ( .A1(n266), .A2(n265), .B1(n263), .B2(n264), .ZN(n262) );
  AOI221D0 U373 ( .A1(n266), .A2(n265), .B1(n264), .B2(n263), .C(n262), .ZN(
        n267) );
  ND4D0 U374 ( .A1(n270), .A2(n269), .A3(n268), .A4(n267), .ZN(n291) );
  NR2D0 U375 ( .A1(n272), .A2(n271), .ZN(n279) );
  MUX2ND0 U376 ( .I0(\DP_OP_13J3_123_8774/n595 ), .I1(n274), .S(n273), .ZN(
        n276) );
  AOI22D0 U377 ( .A1(n279), .A2(n278), .B1(n276), .B2(n277), .ZN(n275) );
  OAI221D0 U378 ( .A1(n279), .A2(n278), .B1(n277), .B2(n276), .C(n275), .ZN(
        n290) );
  CKND2D0 U379 ( .A1(n283), .A2(n282), .ZN(n286) );
  AOI22D0 U380 ( .A1(n287), .A2(n288), .B1(n285), .B2(n286), .ZN(n284) );
  OAI221D0 U381 ( .A1(n288), .A2(n287), .B1(n286), .B2(n285), .C(n284), .ZN(
        n289) );
  NR4D0 U382 ( .A1(n292), .A2(n291), .A3(n290), .A4(n289), .ZN(n302) );
  INVD0 U383 ( .I(\DP_OP_13J3_123_8774/n626 ), .ZN(n294) );
  MUX2ND0 U384 ( .I0(n294), .I1(\DP_OP_13J3_123_8774/n626 ), .S(n293), .ZN(
        n300) );
  CKND2D0 U385 ( .A1(n296), .A2(n295), .ZN(n298) );
  ND3D0 U386 ( .A1(n300), .A2(n299), .A3(n298), .ZN(n297) );
  OAI31D0 U387 ( .A1(n300), .A2(n299), .A3(n298), .B(n297), .ZN(n301) );
  ND4D0 U388 ( .A1(n304), .A2(n303), .A3(n302), .A4(n301), .ZN(n397) );
  NR2D0 U389 ( .A1(n306), .A2(n305), .ZN(n1027) );
  AOI21D0 U390 ( .A1(n1012), .A2(n1027), .B(Q_mag[22]), .ZN(n311) );
  INVD0 U391 ( .I(n311), .ZN(n308) );
  AOI21D0 U392 ( .A1(n1013), .A2(n1027), .B(Q_mag[21]), .ZN(n307) );
  INVD0 U393 ( .I(n307), .ZN(n309) );
  MUX2ND0 U394 ( .I0(n644), .I1(n600), .S(n309), .ZN(n561) );
  NR2D0 U395 ( .A1(n308), .A2(n561), .ZN(n571) );
  AOI33D0 U396 ( .A1(n308), .A2(n600), .A3(n307), .B1(n311), .B2(n644), .B3(
        n309), .ZN(n584) );
  INVD0 U397 ( .I(n584), .ZN(n572) );
  AOI22D0 U398 ( .A1(S_mag[22]), .A2(n571), .B1(S_mag[21]), .B2(n572), .ZN(
        n313) );
  CKND2D0 U399 ( .A1(n644), .A2(n309), .ZN(n310) );
  NR2D0 U400 ( .A1(n311), .A2(n561), .ZN(n570) );
  CKND2D0 U401 ( .A1(n313), .A2(n312), .ZN(n327) );
  AOI21D0 U402 ( .A1(n1023), .A2(n446), .B(Q_mag[19]), .ZN(n314) );
  MUX2ND0 U403 ( .I0(n600), .I1(n644), .S(n314), .ZN(n441) );
  AOI21D0 U404 ( .A1(n1023), .A2(n1012), .B(Q_mag[18]), .ZN(n316) );
  INVD0 U405 ( .I(n316), .ZN(n315) );
  MUX2ND0 U406 ( .I0(n698), .I1(n1029), .S(n315), .ZN(n442) );
  MUX2ND0 U407 ( .I0(n316), .I1(n315), .S(n314), .ZN(n322) );
  IND3D0 U408 ( .A1(n441), .B1(n442), .B2(n322), .ZN(n638) );
  NR2D0 U409 ( .A1(n442), .A2(n441), .ZN(n642) );
  INVD0 U410 ( .I(n642), .ZN(n443) );
  OAI22D0 U411 ( .A1(n933), .A2(n638), .B1(n928), .B2(n443), .ZN(n317) );
  MUX2ND0 U412 ( .I0(n644), .I1(n600), .S(n317), .ZN(n326) );
  INVD0 U413 ( .I(n573), .ZN(n509) );
  INVD0 U414 ( .I(S_mag[19]), .ZN(n850) );
  NR2D0 U415 ( .A1(n509), .A2(n850), .ZN(n319) );
  INVD0 U416 ( .I(n571), .ZN(n585) );
  INVD0 U417 ( .I(S_mag[20]), .ZN(n846) );
  OAI22D0 U418 ( .A1(n930), .A2(n585), .B1(n846), .B2(n584), .ZN(n318) );
  AOI211D0 U419 ( .A1(n941), .A2(n570), .B(n319), .C(n318), .ZN(n325) );
  INVD0 U420 ( .I(S_mag[18]), .ZN(n854) );
  NR2D0 U421 ( .A1(n854), .A2(n509), .ZN(n321) );
  OAI22D0 U422 ( .A1(n846), .A2(n585), .B1(n584), .B2(n850), .ZN(n320) );
  AOI211D0 U423 ( .A1(n945), .A2(n570), .B(n321), .C(n320), .ZN(n337) );
  IND2D0 U424 ( .A1(n322), .B1(n442), .ZN(n639) );
  OAI222D0 U425 ( .A1(n638), .A2(n930), .B1(n639), .B2(n933), .C1(n935), .C2(
        n443), .ZN(n323) );
  MUX2ND0 U426 ( .I0(n644), .I1(n600), .S(n323), .ZN(n336) );
  FA1D0 U427 ( .A(\DP_OP_13J3_123_8774/n477 ), .B(\DP_OP_13J3_123_8774/n470 ), 
        .CI(n324), .CO(n356), .S(n398) );
  NR4D0 U428 ( .A1(\DP_OP_13J3_123_8774/n443 ), .A2(\DP_OP_13J3_123_8774/n460 ), .A3(\DP_OP_13J3_123_8774/n461 ), .A4(n356), .ZN(n364) );
  CKND2D0 U429 ( .A1(n364), .A2(n358), .ZN(n348) );
  NR2D0 U430 ( .A1(\DP_OP_13J3_123_8774/n435 ), .A2(n348), .ZN(n361) );
  INVD0 U431 ( .I(\DP_OP_13J3_123_8774/n423 ), .ZN(n359) );
  CKND2D0 U432 ( .A1(n361), .A2(n359), .ZN(n341) );
  NR2D0 U433 ( .A1(\DP_OP_13J3_123_8774/n417 ), .A2(n341), .ZN(n370) );
  INVD0 U434 ( .I(\DP_OP_13J3_123_8774/n416 ), .ZN(n367) );
  NR2D0 U435 ( .A1(\DP_OP_13J3_123_8774/n406 ), .A2(n365), .ZN(n340) );
  INR2D0 U436 ( .A1(n340), .B1(\DP_OP_13J3_123_8774/n402 ), .ZN(n382) );
  INVD0 U437 ( .I(\DP_OP_13J3_123_8774/n401 ), .ZN(n383) );
  CKAN2D0 U438 ( .A1(n382), .A2(n383), .Z(n329) );
  INR2D0 U439 ( .A1(n329), .B1(\DP_OP_13J3_123_8774/n394 ), .ZN(n380) );
  CKND2D0 U440 ( .A1(n381), .A2(n380), .ZN(n379) );
  INR2D0 U441 ( .A1(n339), .B1(n379), .ZN(n390) );
  INVD0 U442 ( .I(n390), .ZN(n334) );
  FA1D0 U443 ( .A(\DP_OP_13J3_123_8774/n388 ), .B(n326), .CI(n325), .CO(n328), 
        .S(n339) );
  XOR4D0 U444 ( .A1(n600), .A2(\DP_OP_13J3_123_8774/n388 ), .A3(n328), .A4(
        n327), .Z(n333) );
  INVD0 U445 ( .I(\DP_OP_13J3_123_8774/n394 ), .ZN(n330) );
  MUX2ND0 U446 ( .I0(n330), .I1(\DP_OP_13J3_123_8774/n394 ), .S(n329), .ZN(
        n332) );
  NR2D0 U447 ( .A1(n332), .A2(\DP_OP_13J3_123_8774/n396 ), .ZN(n331) );
  AOI221D0 U448 ( .A1(n334), .A2(n333), .B1(\DP_OP_13J3_123_8774/n396 ), .B2(
        n332), .C(n331), .ZN(n335) );
  INVD0 U449 ( .I(n570), .ZN(n587) );
  OA222D0 U450 ( .A1(n933), .A2(n584), .B1(n935), .B2(n587), .C1(n930), .C2(
        n509), .Z(n389) );
  OAI22D0 U451 ( .A1(n933), .A2(n509), .B1(n928), .B2(n587), .ZN(n387) );
  FA1D0 U452 ( .A(\DP_OP_13J3_123_8774/n388 ), .B(n337), .CI(n336), .CO(n338), 
        .S(n381) );
  XNR3D0 U453 ( .A1(n339), .A2(n338), .A3(n379), .ZN(n394) );
  XNR3D0 U454 ( .A1(\DP_OP_13J3_123_8774/n402 ), .A2(n340), .A3(
        \DP_OP_13J3_123_8774/n405 ), .ZN(n378) );
  INVD0 U455 ( .I(n341), .ZN(n347) );
  INVD0 U456 ( .I(\DP_OP_13J3_123_8774/n417 ), .ZN(n342) );
  MUX2ND0 U457 ( .I0(n342), .I1(\DP_OP_13J3_123_8774/n417 ), .S(
        \DP_OP_13J3_123_8774/n422 ), .ZN(n346) );
  INVD0 U458 ( .I(n356), .ZN(n343) );
  MUX2ND0 U459 ( .I0(n356), .I1(n343), .S(\DP_OP_13J3_123_8774/n469 ), .ZN(
        n345) );
  AOI22D0 U460 ( .A1(n347), .A2(n346), .B1(\DP_OP_13J3_123_8774/n461 ), .B2(
        n345), .ZN(n344) );
  OAI221D0 U461 ( .A1(n347), .A2(n346), .B1(n345), .B2(
        \DP_OP_13J3_123_8774/n461 ), .C(n344), .ZN(n377) );
  MUX2ND0 U462 ( .I0(n349), .I1(\DP_OP_13J3_123_8774/n435 ), .S(
        \DP_OP_13J3_123_8774/n428 ), .ZN(n354) );
  NR3D0 U463 ( .A1(\DP_OP_13J3_123_8774/n460 ), .A2(\DP_OP_13J3_123_8774/n461 ), .A3(n356), .ZN(n353) );
  INVD0 U464 ( .I(\DP_OP_13J3_123_8774/n443 ), .ZN(n350) );
  MUX2ND0 U465 ( .I0(n350), .I1(\DP_OP_13J3_123_8774/n443 ), .S(
        \DP_OP_13J3_123_8774/n450 ), .ZN(n352) );
  AOI22D0 U466 ( .A1(n355), .A2(n354), .B1(n353), .B2(n352), .ZN(n351) );
  OAI221D0 U467 ( .A1(n355), .A2(n354), .B1(n353), .B2(n352), .C(n351), .ZN(
        n376) );
  NR2D0 U468 ( .A1(\DP_OP_13J3_123_8774/n461 ), .A2(n356), .ZN(n357) );
  XOR3D0 U469 ( .A1(\DP_OP_13J3_123_8774/n460 ), .A2(n357), .A3(
        \DP_OP_13J3_123_8774/n451 ), .Z(n374) );
  MUX2ND0 U470 ( .I0(n358), .I1(\DP_OP_13J3_123_8774/n436 ), .S(
        \DP_OP_13J3_123_8774/n442 ), .ZN(n363) );
  MUX2ND0 U471 ( .I0(n359), .I1(\DP_OP_13J3_123_8774/n423 ), .S(
        \DP_OP_13J3_123_8774/n427 ), .ZN(n362) );
  OAI22D0 U472 ( .A1(n364), .A2(n363), .B1(n361), .B2(n362), .ZN(n360) );
  AOI221D0 U473 ( .A1(n364), .A2(n363), .B1(n362), .B2(n361), .C(n360), .ZN(
        n373) );
  INVD0 U474 ( .I(\DP_OP_13J3_123_8774/n406 ), .ZN(n366) );
  MUX2ND0 U475 ( .I0(\DP_OP_13J3_123_8774/n406 ), .I1(n366), .S(n365), .ZN(
        n371) );
  MUX2ND0 U476 ( .I0(n367), .I1(\DP_OP_13J3_123_8774/n416 ), .S(
        \DP_OP_13J3_123_8774/n410 ), .ZN(n369) );
  OAI22D0 U477 ( .A1(\DP_OP_13J3_123_8774/n409 ), .A2(n371), .B1(n370), .B2(
        n369), .ZN(n368) );
  AOI221D0 U478 ( .A1(n371), .A2(\DP_OP_13J3_123_8774/n409 ), .B1(n370), .B2(
        n369), .C(n368), .ZN(n372) );
  ND4D0 U479 ( .A1(running), .A2(n374), .A3(n373), .A4(n372), .ZN(n375) );
  NR4D0 U480 ( .A1(n378), .A2(n377), .A3(n376), .A4(n375), .ZN(n393) );
  MUX2ND0 U481 ( .I0(n383), .I1(\DP_OP_13J3_123_8774/n401 ), .S(n382), .ZN(
        n385) );
  OAI22D0 U482 ( .A1(\DP_OP_13J3_123_8774/n397 ), .A2(n385), .B1(
        \DP_OP_13J3_123_8774/n393 ), .B2(n386), .ZN(n384) );
  AOI221D0 U483 ( .A1(n386), .A2(\DP_OP_13J3_123_8774/n393 ), .B1(n385), .B2(
        \DP_OP_13J3_123_8774/n397 ), .C(n384), .ZN(n392) );
  OAI31D0 U484 ( .A1(n390), .A2(n389), .A3(n388), .B(n387), .ZN(n391) );
  ND4D0 U485 ( .A1(n394), .A2(n393), .A3(n392), .A4(n391), .ZN(n395) );
  AO211D0 U486 ( .A1(n398), .A2(n397), .B(n396), .C(n395), .Z(n1016) );
  OAI22D0 U487 ( .A1(n400), .A2(n399), .B1(n405), .B2(n1016), .ZN(n67) );
  NR2D0 U488 ( .A1(n405), .A2(n404), .ZN(N67) );
  CKND2D0 U489 ( .A1(n1025), .A2(n1011), .ZN(n72) );
  NR3D0 U490 ( .A1(bit_pos[4]), .A2(n407), .A3(n406), .ZN(n1020) );
  AOI21D0 U491 ( .A1(n1020), .A2(n1017), .B(Q_mag[12]), .ZN(n410) );
  INVD0 U492 ( .I(n410), .ZN(n409) );
  MUX2ND0 U493 ( .I0(n828), .I1(n1030), .S(n409), .ZN(n412) );
  NR2D0 U494 ( .A1(n583), .A2(n412), .ZN(n568) );
  AOI21D0 U495 ( .A1(n1020), .A2(n1013), .B(Q_mag[13]), .ZN(n408) );
  MUX2ND0 U496 ( .I0(n709), .I1(n774), .S(n408), .ZN(n413) );
  NR2D0 U497 ( .A1(n412), .A2(n413), .ZN(n772) );
  INVD0 U498 ( .I(n772), .ZN(n707) );
  IND2D0 U499 ( .A1(n412), .B1(n413), .ZN(n768) );
  MUX2ND0 U500 ( .I0(n410), .I1(n409), .S(n408), .ZN(n411) );
  IND2D0 U501 ( .A1(n411), .B1(n412), .ZN(n767) );
  OAI222D0 U502 ( .A1(n707), .A2(n586), .B1(n768), .B2(n921), .C1(n767), .C2(
        n583), .ZN(n435) );
  INVD0 U503 ( .I(n435), .ZN(n436) );
  IND3D0 U504 ( .A1(n568), .B1(n774), .B2(n436), .ZN(n417) );
  NR2D0 U505 ( .A1(n921), .A2(n767), .ZN(n415) );
  IND3D0 U506 ( .A1(n413), .B1(n412), .B2(n411), .ZN(n769) );
  OAI22D0 U507 ( .A1(n917), .A2(n768), .B1(n583), .B2(n769), .ZN(n414) );
  AOI211D0 U508 ( .A1(n772), .A2(n542), .B(n415), .C(n414), .ZN(n418) );
  CKND2D0 U509 ( .A1(n418), .A2(n774), .ZN(n416) );
  NR2D0 U510 ( .A1(n417), .A2(n416), .ZN(\DP_OP_13J3_123_8774/n598 ) );
  MUX2ND0 U511 ( .I0(n927), .I1(n839), .S(n420), .ZN(n423) );
  INVD0 U512 ( .I(n423), .ZN(n424) );
  NR2D0 U513 ( .A1(n583), .A2(n424), .ZN(\DP_OP_13J3_123_8774/n628 ) );
  OAI211D0 U514 ( .A1(n418), .A2(n774), .B(n417), .C(n416), .ZN(n419) );
  IND2D0 U515 ( .A1(\DP_OP_13J3_123_8774/n598 ), .B1(n419), .ZN(n559) );
  AOI21D0 U516 ( .A1(n1019), .A2(n1012), .B(Q_mag[10]), .ZN(n421) );
  XNR2D0 U517 ( .A1(n420), .A2(n421), .ZN(n422) );
  MUX2ND0 U518 ( .I0(n828), .I1(n1030), .S(n421), .ZN(n425) );
  ND3D0 U519 ( .A1(n424), .A2(n422), .A3(n425), .ZN(n778) );
  INVD0 U520 ( .I(n778), .ZN(n830) );
  CKND2D0 U521 ( .A1(n423), .A2(n425), .ZN(n776) );
  INVD0 U522 ( .I(n776), .ZN(n829) );
  AOI22D0 U523 ( .A1(S_mag[2]), .A2(n830), .B1(n914), .B2(n829), .ZN(n427) );
  NR2D0 U524 ( .A1(n423), .A2(n422), .ZN(n832) );
  NR2D0 U525 ( .A1(n425), .A2(n424), .ZN(n831) );
  AOI22D0 U526 ( .A1(S_mag[3]), .A2(n832), .B1(S_mag[4]), .B2(n831), .ZN(n426)
         );
  CKND2D0 U527 ( .A1(n427), .A2(n426), .ZN(n428) );
  MUX2ND0 U528 ( .I0(n828), .I1(n1030), .S(n428), .ZN(n555) );
  AOI22D0 U529 ( .A1(S_mag[0]), .A2(n830), .B1(n542), .B2(n829), .ZN(n430) );
  AOI22D0 U530 ( .A1(S_mag[2]), .A2(n831), .B1(S_mag[1]), .B2(n832), .ZN(n429)
         );
  CKND2D0 U531 ( .A1(n430), .A2(n429), .ZN(n551) );
  NR2D0 U532 ( .A1(n1030), .A2(n551), .ZN(n550) );
  AOI222D0 U533 ( .A1(n829), .A2(n462), .B1(n831), .B2(S_mag[1]), .C1(n832), 
        .C2(S_mag[0]), .ZN(n581) );
  INVD0 U534 ( .I(n581), .ZN(n582) );
  NR3D0 U535 ( .A1(n1030), .A2(\DP_OP_13J3_123_8774/n628 ), .A3(n582), .ZN(
        n549) );
  CKAN2D0 U536 ( .A1(n550), .A2(n549), .Z(n566) );
  AOI22D0 U537 ( .A1(S_mag[1]), .A2(n830), .B1(n924), .B2(n829), .ZN(n432) );
  AOI22D0 U538 ( .A1(S_mag[2]), .A2(n832), .B1(S_mag[3]), .B2(n831), .ZN(n431)
         );
  CKND2D0 U539 ( .A1(n432), .A2(n431), .ZN(n433) );
  MUX2ND0 U540 ( .I0(n1030), .I1(n828), .S(n433), .ZN(n567) );
  OAI21D0 U541 ( .A1(n566), .A2(n568), .B(n567), .ZN(n554) );
  CKND2D0 U542 ( .A1(n568), .A2(n774), .ZN(n434) );
  MUX2ND0 U543 ( .I0(n436), .I1(n435), .S(n434), .ZN(n553) );
  AOI22D0 U544 ( .A1(S_mag[3]), .A2(n830), .B1(n909), .B2(n829), .ZN(n438) );
  AOI22D0 U545 ( .A1(S_mag[4]), .A2(n832), .B1(S_mag[5]), .B2(n831), .ZN(n437)
         );
  CKND2D0 U546 ( .A1(n438), .A2(n437), .ZN(n439) );
  MUX2ND0 U547 ( .I0(n828), .I1(n1030), .S(n439), .ZN(n557) );
  INVD0 U548 ( .I(n440), .ZN(\DP_OP_13J3_123_8774/n596 ) );
  NR2D0 U549 ( .A1(n583), .A2(n442), .ZN(n565) );
  IND2D0 U550 ( .A1(n442), .B1(n441), .ZN(n637) );
  OAI222D0 U551 ( .A1(n443), .A2(n586), .B1(n637), .B2(n921), .C1(n583), .C2(
        n639), .ZN(n467) );
  INVD0 U552 ( .I(n467), .ZN(n468) );
  IND3D0 U553 ( .A1(n565), .B1(n644), .B2(n468), .ZN(n448) );
  NR2D0 U554 ( .A1(n917), .A2(n637), .ZN(n445) );
  OAI22D0 U555 ( .A1(n921), .A2(n639), .B1(n583), .B2(n638), .ZN(n444) );
  AOI211D0 U556 ( .A1(n642), .A2(n542), .B(n445), .C(n444), .ZN(n449) );
  CKND2D0 U557 ( .A1(n449), .A2(n644), .ZN(n447) );
  NR2D0 U558 ( .A1(n448), .A2(n447), .ZN(\DP_OP_13J3_123_8774/n547 ) );
  MUX2ND0 U559 ( .I0(n774), .I1(n709), .S(n451), .ZN(n454) );
  INVD0 U560 ( .I(n454), .ZN(n455) );
  NR2D0 U561 ( .A1(n583), .A2(n455), .ZN(\DP_OP_13J3_123_8774/n592 ) );
  OAI211D0 U562 ( .A1(n449), .A2(n644), .B(n448), .C(n447), .ZN(n450) );
  IND2D0 U563 ( .A1(\DP_OP_13J3_123_8774/n547 ), .B1(n450), .ZN(n547) );
  AOI21D0 U564 ( .A1(n1023), .A2(n1017), .B(Q_mag[16]), .ZN(n452) );
  XNR2D0 U565 ( .A1(n451), .A2(n452), .ZN(n453) );
  MUX2ND0 U566 ( .I0(n698), .I1(n1029), .S(n452), .ZN(n456) );
  ND3D0 U567 ( .A1(n455), .A2(n453), .A3(n456), .ZN(n648) );
  INVD0 U568 ( .I(n648), .ZN(n700) );
  CKND2D0 U569 ( .A1(n454), .A2(n456), .ZN(n646) );
  AOI22D0 U570 ( .A1(S_mag[2]), .A2(n700), .B1(n914), .B2(n699), .ZN(n458) );
  NR2D0 U571 ( .A1(n454), .A2(n453), .ZN(n702) );
  NR2D0 U572 ( .A1(n456), .A2(n455), .ZN(n701) );
  CKND2D0 U573 ( .A1(n458), .A2(n457), .ZN(n459) );
  MUX2ND0 U574 ( .I0(n698), .I1(n1029), .S(n459), .ZN(n540) );
  AOI22D0 U575 ( .A1(S_mag[0]), .A2(n700), .B1(n542), .B2(n699), .ZN(n461) );
  AOI22D0 U576 ( .A1(S_mag[2]), .A2(n701), .B1(S_mag[1]), .B2(n702), .ZN(n460)
         );
  CKND2D0 U577 ( .A1(n461), .A2(n460), .ZN(n536) );
  NR2D0 U578 ( .A1(n1029), .A2(n536), .ZN(n535) );
  AOI222D0 U579 ( .A1(n699), .A2(n462), .B1(n701), .B2(S_mag[1]), .C1(n702), 
        .C2(S_mag[0]), .ZN(n578) );
  INVD0 U580 ( .I(n578), .ZN(n579) );
  NR3D0 U581 ( .A1(n1029), .A2(\DP_OP_13J3_123_8774/n592 ), .A3(n579), .ZN(
        n534) );
  CKAN2D0 U582 ( .A1(n535), .A2(n534), .Z(n563) );
  AOI22D0 U583 ( .A1(S_mag[1]), .A2(n700), .B1(n924), .B2(n699), .ZN(n464) );
  AOI22D0 U584 ( .A1(S_mag[2]), .A2(n702), .B1(S_mag[3]), .B2(n701), .ZN(n463)
         );
  CKND2D0 U585 ( .A1(n464), .A2(n463), .ZN(n465) );
  MUX2ND0 U586 ( .I0(n1029), .I1(n698), .S(n465), .ZN(n564) );
  OAI21D0 U587 ( .A1(n563), .A2(n565), .B(n564), .ZN(n539) );
  CKND2D0 U588 ( .A1(n565), .A2(n644), .ZN(n466) );
  MUX2ND0 U589 ( .I0(n468), .I1(n467), .S(n466), .ZN(n538) );
  AOI22D0 U590 ( .A1(S_mag[3]), .A2(n700), .B1(n909), .B2(n699), .ZN(n470) );
  AOI22D0 U591 ( .A1(S_mag[4]), .A2(n702), .B1(S_mag[5]), .B2(n701), .ZN(n469)
         );
  CKND2D0 U592 ( .A1(n470), .A2(n469), .ZN(n471) );
  MUX2ND0 U593 ( .I0(n698), .I1(n1029), .S(n471), .ZN(n545) );
  INVD0 U594 ( .I(n472), .ZN(\DP_OP_13J3_123_8774/n545 ) );
  FA1D0 U595 ( .A(n475), .B(n474), .CI(n473), .CO(n476), .S(n296) );
  INVD0 U596 ( .I(n476), .ZN(\DP_OP_13J3_123_8774/n629 ) );
  AOI22D0 U597 ( .A1(S_mag[13]), .A2(n571), .B1(n973), .B2(n570), .ZN(n478) );
  AOI22D0 U598 ( .A1(S_mag[12]), .A2(n572), .B1(S_mag[11]), .B2(n573), .ZN(
        n477) );
  CKND2D0 U599 ( .A1(n478), .A2(n477), .ZN(\DP_OP_13J3_123_8774/n727 ) );
  AOI22D0 U600 ( .A1(S_mag[7]), .A2(n571), .B1(n997), .B2(n570), .ZN(n480) );
  AOI22D0 U601 ( .A1(S_mag[5]), .A2(n573), .B1(S_mag[6]), .B2(n572), .ZN(n479)
         );
  CKND2D0 U602 ( .A1(n480), .A2(n479), .ZN(\DP_OP_13J3_123_8774/n732 ) );
  AOI22D0 U603 ( .A1(S_mag[18]), .A2(n572), .B1(n571), .B2(S_mag[19]), .ZN(
        n482) );
  AOI22D0 U604 ( .A1(S_mag[17]), .A2(n573), .B1(n570), .B2(n949), .ZN(n481) );
  CKND2D0 U605 ( .A1(n482), .A2(n481), .ZN(\DP_OP_13J3_123_8774/n721 ) );
  INVD0 U606 ( .I(S_mag[17]), .ZN(n858) );
  NR2D0 U607 ( .A1(n858), .A2(n637), .ZN(n484) );
  INVD0 U608 ( .I(S_mag[15]), .ZN(n866) );
  INVD0 U609 ( .I(S_mag[16]), .ZN(n862) );
  OAI22D0 U610 ( .A1(n866), .A2(n638), .B1(n862), .B2(n639), .ZN(n483) );
  AOI211D0 U611 ( .A1(n642), .A2(n957), .B(n484), .C(n483), .ZN(n485) );
  MUX2ND0 U612 ( .I0(n600), .I1(n644), .S(n485), .ZN(n518) );
  INVD0 U613 ( .I(S_mag[12]), .ZN(n878) );
  NR2D0 U614 ( .A1(n878), .A2(n509), .ZN(n487) );
  INVD0 U615 ( .I(S_mag[14]), .ZN(n870) );
  INVD0 U616 ( .I(S_mag[13]), .ZN(n874) );
  OAI22D0 U617 ( .A1(n870), .A2(n585), .B1(n874), .B2(n584), .ZN(n486) );
  AOI211D0 U618 ( .A1(n570), .A2(n969), .B(n487), .C(n486), .ZN(n517) );
  NR2D0 U619 ( .A1(n874), .A2(n509), .ZN(n489) );
  AOI211D0 U620 ( .A1(n570), .A2(n965), .B(n489), .C(n488), .ZN(n501) );
  INVD0 U621 ( .I(n490), .ZN(\DP_OP_13J3_123_8774/n411 ) );
  AOI22D0 U622 ( .A1(S_mag[5]), .A2(n571), .B1(n909), .B2(n570), .ZN(n492) );
  AOI22D0 U623 ( .A1(S_mag[3]), .A2(n573), .B1(S_mag[4]), .B2(n572), .ZN(n491)
         );
  CKND2D0 U624 ( .A1(n492), .A2(n491), .ZN(\DP_OP_13J3_123_8774/n734 ) );
  INVD0 U625 ( .I(S_mag[11]), .ZN(n882) );
  NR2D0 U626 ( .A1(n882), .A2(n637), .ZN(n494) );
  INVD0 U627 ( .I(S_mag[9]), .ZN(n890) );
  INVD0 U628 ( .I(S_mag[10]), .ZN(n886) );
  OAI22D0 U629 ( .A1(n890), .A2(n638), .B1(n886), .B2(n639), .ZN(n493) );
  MUX2ND0 U630 ( .I0(n600), .I1(n644), .S(n495), .ZN(n530) );
  INVD0 U631 ( .I(S_mag[6]), .ZN(n902) );
  NR2D0 U632 ( .A1(n902), .A2(n509), .ZN(n497) );
  INVD0 U633 ( .I(S_mag[7]), .ZN(n898) );
  INVD0 U634 ( .I(S_mag[8]), .ZN(n894) );
  OAI22D0 U635 ( .A1(n898), .A2(n584), .B1(n894), .B2(n585), .ZN(n496) );
  AOI211D0 U636 ( .A1(n570), .A2(n993), .B(n497), .C(n496), .ZN(n529) );
  AOI22D0 U637 ( .A1(S_mag[4]), .A2(n571), .B1(n914), .B2(n570), .ZN(n500) );
  AOI22D0 U638 ( .A1(S_mag[2]), .A2(n573), .B1(S_mag[3]), .B2(n572), .ZN(n499)
         );
  CKND2D0 U639 ( .A1(n500), .A2(n499), .ZN(\DP_OP_13J3_123_8774/n735 ) );
  FA1D0 U640 ( .A(\DP_OP_13J3_123_8774/n413 ), .B(n502), .CI(n501), .CO(n490), 
        .S(n503) );
  INVD0 U641 ( .I(n503), .ZN(\DP_OP_13J3_123_8774/n412 ) );
  AOI22D0 U642 ( .A1(S_mag[12]), .A2(n571), .B1(n977), .B2(n570), .ZN(n505) );
  AOI22D0 U643 ( .A1(S_mag[10]), .A2(n573), .B1(S_mag[11]), .B2(n572), .ZN(
        n504) );
  CKND2D0 U644 ( .A1(n505), .A2(n504), .ZN(\DP_OP_13J3_123_8774/n728 ) );
  NR2D0 U645 ( .A1(n882), .A2(n639), .ZN(n507) );
  OAI22D0 U646 ( .A1(n886), .A2(n638), .B1(n878), .B2(n637), .ZN(n506) );
  AOI211D0 U647 ( .A1(n642), .A2(n977), .B(n507), .C(n506), .ZN(n508) );
  MUX2ND0 U648 ( .I0(n600), .I1(n644), .S(n508), .ZN(n521) );
  NR2D0 U649 ( .A1(n898), .A2(n509), .ZN(n511) );
  OAI22D0 U650 ( .A1(n894), .A2(n584), .B1(n890), .B2(n585), .ZN(n510) );
  AOI211D0 U651 ( .A1(n570), .A2(n989), .B(n511), .C(n510), .ZN(n520) );
  INVD0 U652 ( .I(n512), .ZN(\DP_OP_13J3_123_8774/n456 ) );
  AOI22D0 U653 ( .A1(S_mag[6]), .A2(n571), .B1(n1002), .B2(n570), .ZN(n514) );
  AOI22D0 U654 ( .A1(S_mag[4]), .A2(n573), .B1(S_mag[5]), .B2(n572), .ZN(n513)
         );
  AOI22D0 U655 ( .A1(S_mag[17]), .A2(n572), .B1(S_mag[18]), .B2(n571), .ZN(
        n516) );
  AOI22D0 U656 ( .A1(S_mag[16]), .A2(n573), .B1(n953), .B2(n570), .ZN(n515) );
  CKND2D0 U657 ( .A1(n516), .A2(n515), .ZN(\DP_OP_13J3_123_8774/n722 ) );
  FA1D0 U658 ( .A(\DP_OP_13J3_123_8774/n413 ), .B(n518), .CI(n517), .CO(n502), 
        .S(n519) );
  INVD0 U659 ( .I(n519), .ZN(\DP_OP_13J3_123_8774/n419 ) );
  FA1D0 U660 ( .A(\DP_OP_13J3_123_8774/n457 ), .B(n521), .CI(n520), .CO(n522), 
        .S(n512) );
  INVD0 U661 ( .I(n522), .ZN(\DP_OP_13J3_123_8774/n455 ) );
  AOI22D0 U662 ( .A1(S_mag[16]), .A2(n571), .B1(n570), .B2(n961), .ZN(n524) );
  AOI22D0 U663 ( .A1(S_mag[14]), .A2(n573), .B1(S_mag[15]), .B2(n572), .ZN(
        n523) );
  CKND2D0 U664 ( .A1(n524), .A2(n523), .ZN(n569) );
  INVD0 U665 ( .I(\DP_OP_13J3_123_8774/n398 ), .ZN(\DP_OP_13J3_123_8774/n403 )
         );
  AOI22D0 U666 ( .A1(S_mag[3]), .A2(n571), .B1(n924), .B2(n570), .ZN(n526) );
  AOI22D0 U667 ( .A1(S_mag[2]), .A2(n572), .B1(S_mag[1]), .B2(n573), .ZN(n525)
         );
  AOI22D0 U668 ( .A1(S_mag[17]), .A2(n571), .B1(S_mag[16]), .B2(n572), .ZN(
        n528) );
  AOI22D0 U669 ( .A1(S_mag[15]), .A2(n573), .B1(n957), .B2(n570), .ZN(n527) );
  FA1D0 U670 ( .A(\DP_OP_13J3_123_8774/n457 ), .B(n530), .CI(n529), .CO(n531), 
        .S(n498) );
  INVD0 U671 ( .I(n531), .ZN(\DP_OP_13J3_123_8774/n465 ) );
  AOI22D0 U672 ( .A1(S_mag[9]), .A2(n573), .B1(S_mag[10]), .B2(n572), .ZN(n532) );
  CKND2D0 U673 ( .A1(n533), .A2(n532), .ZN(\DP_OP_13J3_123_8774/n432 ) );
  INVD0 U674 ( .I(\DP_OP_13J3_123_8774/n432 ), .ZN(\DP_OP_13J3_123_8774/n440 )
         );
  AOI211D0 U675 ( .A1(n1029), .A2(n536), .B(n535), .C(n534), .ZN(n537) );
  NR2D0 U676 ( .A1(n563), .A2(n537), .ZN(\DP_OP_13J3_123_8774/n576 ) );
  FA1D0 U677 ( .A(n540), .B(n539), .CI(n538), .CO(n546), .S(n541) );
  INVD0 U678 ( .I(n541), .ZN(\DP_OP_13J3_123_8774/n556 ) );
  AOI22D0 U679 ( .A1(S_mag[2]), .A2(n571), .B1(n542), .B2(n570), .ZN(n544) );
  AOI22D0 U680 ( .A1(S_mag[1]), .A2(n572), .B1(S_mag[0]), .B2(n573), .ZN(n543)
         );
  FA1D0 U681 ( .A(n547), .B(n546), .CI(n545), .CO(n472), .S(n548) );
  AOI211D0 U682 ( .A1(n1030), .A2(n551), .B(n550), .C(n549), .ZN(n552) );
  NR2D0 U683 ( .A1(n566), .A2(n552), .ZN(\DP_OP_13J3_123_8774/n618 ) );
  FA1D0 U684 ( .A(n555), .B(n554), .CI(n553), .CO(n558), .S(n556) );
  INVD0 U685 ( .I(n556), .ZN(\DP_OP_13J3_123_8774/n604 ) );
  FA1D0 U686 ( .A(n559), .B(n558), .CI(n557), .CO(n440), .S(n560) );
  INVD0 U687 ( .I(n560), .ZN(\DP_OP_13J3_123_8774/n597 ) );
  NR2D0 U688 ( .A1(n583), .A2(n561), .ZN(\DP_OP_13J3_123_8774/n739 ) );
  IOA21D0 U689 ( .A1(bit_pos[4]), .A2(n562), .B(n1025), .ZN(n73) );
  XOR3D0 U690 ( .A1(n565), .A2(n564), .A3(n563), .Z(\DP_OP_13J3_123_8774/n566 ) );
  XOR3D0 U691 ( .A1(n568), .A2(n567), .A3(n566), .Z(\DP_OP_13J3_123_8774/n611 ) );
  FA1D0 U692 ( .A(\DP_OP_13J3_123_8774/n413 ), .B(n709), .CI(n569), .CO(
        \DP_OP_13J3_123_8774/n398 ), .S(\DP_OP_13J3_123_8774/n407 ) );
  AOI22D0 U693 ( .A1(S_mag[10]), .A2(n571), .B1(n985), .B2(n570), .ZN(n575) );
  AOI22D0 U694 ( .A1(S_mag[8]), .A2(n573), .B1(S_mag[9]), .B2(n572), .ZN(n574)
         );
  CKND2D0 U695 ( .A1(n575), .A2(n574), .ZN(n576) );
  FA1D0 U696 ( .A(\DP_OP_13J3_123_8774/n457 ), .B(n839), .CI(n576), .CO(
        \DP_OP_13J3_123_8774/n447 ), .S(\DP_OP_13J3_123_8774/n448 ) );
  CKND2D0 U697 ( .A1(\DP_OP_13J3_123_8774/n592 ), .A2(n698), .ZN(n577) );
  MUX2ND0 U698 ( .I0(n579), .I1(n578), .S(n577), .ZN(
        \DP_OP_13J3_123_8774/n584 ) );
  CKND2D0 U699 ( .A1(\DP_OP_13J3_123_8774/n628 ), .A2(n828), .ZN(n580) );
  MUX2ND0 U700 ( .I0(n582), .I1(n581), .S(n580), .ZN(
        \DP_OP_13J3_123_8774/n623 ) );
  OAI222D0 U701 ( .A1(n587), .A2(n586), .B1(n585), .B2(n921), .C1(n584), .C2(
        n583), .ZN(\DP_OP_13J3_123_8774/n738 ) );
  NR2D0 U702 ( .A1(n933), .A2(n637), .ZN(n589) );
  OAI22D0 U703 ( .A1(n930), .A2(n639), .B1(n846), .B2(n638), .ZN(n588) );
  AOI211D0 U704 ( .A1(n642), .A2(n937), .B(n589), .C(n588), .ZN(n590) );
  MUX2ND0 U705 ( .I0(n644), .I1(n600), .S(n590), .ZN(
        \DP_OP_13J3_123_8774/n743 ) );
  NR2D0 U706 ( .A1(n930), .A2(n637), .ZN(n592) );
  OAI22D0 U707 ( .A1(n846), .A2(n639), .B1(n638), .B2(n850), .ZN(n591) );
  AOI211D0 U708 ( .A1(n642), .A2(n941), .B(n592), .C(n591), .ZN(n593) );
  MUX2ND0 U709 ( .I0(n644), .I1(n600), .S(n593), .ZN(
        \DP_OP_13J3_123_8774/n744 ) );
  NR2D0 U710 ( .A1(n846), .A2(n637), .ZN(n595) );
  OAI22D0 U711 ( .A1(n854), .A2(n638), .B1(n639), .B2(n850), .ZN(n594) );
  AOI211D0 U712 ( .A1(n642), .A2(n945), .B(n595), .C(n594), .ZN(n596) );
  MUX2ND0 U713 ( .I0(n644), .I1(n600), .S(n596), .ZN(
        \DP_OP_13J3_123_8774/n745 ) );
  NR2D0 U714 ( .A1(n637), .A2(n850), .ZN(n598) );
  OAI22D0 U715 ( .A1(n858), .A2(n638), .B1(n854), .B2(n639), .ZN(n597) );
  AOI211D0 U716 ( .A1(n642), .A2(n949), .B(n598), .C(n597), .ZN(n599) );
  MUX2ND0 U717 ( .I0(n644), .I1(n600), .S(n599), .ZN(
        \DP_OP_13J3_123_8774/n746 ) );
  NR2D0 U718 ( .A1(n854), .A2(n637), .ZN(n602) );
  OAI22D0 U719 ( .A1(n858), .A2(n639), .B1(n862), .B2(n638), .ZN(n601) );
  AOI211D0 U720 ( .A1(n642), .A2(n953), .B(n602), .C(n601), .ZN(n603) );
  MUX2ND0 U721 ( .I0(n644), .I1(n600), .S(n603), .ZN(
        \DP_OP_13J3_123_8774/n747 ) );
  NR2D0 U722 ( .A1(n862), .A2(n637), .ZN(n605) );
  OAI22D0 U723 ( .A1(n870), .A2(n638), .B1(n866), .B2(n639), .ZN(n604) );
  AOI211D0 U724 ( .A1(n642), .A2(n961), .B(n605), .C(n604), .ZN(n606) );
  MUX2ND0 U725 ( .I0(n644), .I1(n600), .S(n606), .ZN(
        \DP_OP_13J3_123_8774/n749 ) );
  NR2D0 U726 ( .A1(n866), .A2(n637), .ZN(n608) );
  OAI22D0 U727 ( .A1(n870), .A2(n639), .B1(n874), .B2(n638), .ZN(n607) );
  AOI211D0 U728 ( .A1(n642), .A2(n965), .B(n608), .C(n607), .ZN(n609) );
  MUX2ND0 U729 ( .I0(n644), .I1(n600), .S(n609), .ZN(
        \DP_OP_13J3_123_8774/n750 ) );
  NR2D0 U730 ( .A1(n870), .A2(n637), .ZN(n611) );
  OAI22D0 U731 ( .A1(n874), .A2(n639), .B1(n878), .B2(n638), .ZN(n610) );
  AOI211D0 U732 ( .A1(n642), .A2(n969), .B(n611), .C(n610), .ZN(n612) );
  MUX2ND0 U733 ( .I0(n644), .I1(n600), .S(n612), .ZN(
        \DP_OP_13J3_123_8774/n751 ) );
  NR2D0 U734 ( .A1(n878), .A2(n639), .ZN(n614) );
  OAI22D0 U735 ( .A1(n874), .A2(n637), .B1(n882), .B2(n638), .ZN(n613) );
  AOI211D0 U736 ( .A1(n642), .A2(n973), .B(n614), .C(n613), .ZN(n615) );
  MUX2ND0 U737 ( .I0(n644), .I1(n600), .S(n615), .ZN(
        \DP_OP_13J3_123_8774/n752 ) );
  NR2D0 U738 ( .A1(n886), .A2(n637), .ZN(n617) );
  OAI22D0 U739 ( .A1(n894), .A2(n638), .B1(n890), .B2(n639), .ZN(n616) );
  MUX2ND0 U740 ( .I0(n644), .I1(n600), .S(n618), .ZN(
        \DP_OP_13J3_123_8774/n755 ) );
  NR2D0 U741 ( .A1(n890), .A2(n637), .ZN(n620) );
  OAI22D0 U742 ( .A1(n898), .A2(n638), .B1(n894), .B2(n639), .ZN(n619) );
  AOI211D0 U743 ( .A1(n642), .A2(n989), .B(n620), .C(n619), .ZN(n621) );
  MUX2ND0 U744 ( .I0(n644), .I1(n600), .S(n621), .ZN(
        \DP_OP_13J3_123_8774/n756 ) );
  NR2D0 U745 ( .A1(n894), .A2(n637), .ZN(n623) );
  OAI22D0 U746 ( .A1(n902), .A2(n638), .B1(n898), .B2(n639), .ZN(n622) );
  AOI211D0 U747 ( .A1(n642), .A2(n993), .B(n623), .C(n622), .ZN(n624) );
  MUX2ND0 U748 ( .I0(n644), .I1(n600), .S(n624), .ZN(
        \DP_OP_13J3_123_8774/n757 ) );
  NR2D0 U749 ( .A1(n898), .A2(n637), .ZN(n626) );
  INVD0 U750 ( .I(S_mag[5]), .ZN(n906) );
  OAI22D0 U751 ( .A1(n906), .A2(n638), .B1(n902), .B2(n639), .ZN(n625) );
  AOI211D0 U752 ( .A1(n642), .A2(n997), .B(n626), .C(n625), .ZN(n627) );
  MUX2ND0 U753 ( .I0(n644), .I1(n600), .S(n627), .ZN(
        \DP_OP_13J3_123_8774/n758 ) );
  NR2D0 U754 ( .A1(n902), .A2(n637), .ZN(n629) );
  INVD0 U755 ( .I(S_mag[4]), .ZN(n911) );
  AOI211D0 U756 ( .A1(n642), .A2(n1002), .B(n629), .C(n628), .ZN(n630) );
  MUX2ND0 U757 ( .I0(n644), .I1(n600), .S(n630), .ZN(
        \DP_OP_13J3_123_8774/n759 ) );
  NR2D0 U758 ( .A1(n906), .A2(n637), .ZN(n632) );
  INVD0 U759 ( .I(S_mag[3]), .ZN(n919) );
  OAI22D0 U760 ( .A1(n919), .A2(n638), .B1(n911), .B2(n639), .ZN(n631) );
  AOI211D0 U761 ( .A1(n642), .A2(n909), .B(n632), .C(n631), .ZN(n633) );
  MUX2ND0 U762 ( .I0(n644), .I1(n600), .S(n633), .ZN(
        \DP_OP_13J3_123_8774/n760 ) );
  NR2D0 U763 ( .A1(n911), .A2(n637), .ZN(n635) );
  AOI211D0 U764 ( .A1(n642), .A2(n914), .B(n635), .C(n634), .ZN(n636) );
  MUX2ND0 U765 ( .I0(n644), .I1(n600), .S(n636), .ZN(
        \DP_OP_13J3_123_8774/n761 ) );
  OAI22D0 U766 ( .A1(n917), .A2(n639), .B1(n921), .B2(n638), .ZN(n640) );
  AOI211D0 U767 ( .A1(n642), .A2(n924), .B(n641), .C(n640), .ZN(n643) );
  MUX2ND0 U768 ( .I0(n644), .I1(n600), .S(n643), .ZN(
        \DP_OP_13J3_123_8774/n762 ) );
  OAI22D0 U769 ( .A1(n933), .A2(n648), .B1(n928), .B2(n646), .ZN(n645) );
  MUX2ND0 U770 ( .I0(n1029), .I1(n698), .S(n645), .ZN(
        \DP_OP_13J3_123_8774/n767 ) );
  INVD0 U771 ( .I(n702), .ZN(n647) );
  OAI222D0 U772 ( .A1(n648), .A2(n930), .B1(n647), .B2(n933), .C1(n935), .C2(
        n646), .ZN(n649) );
  MUX2ND0 U773 ( .I0(n1029), .I1(n698), .S(n649), .ZN(
        \DP_OP_13J3_123_8774/n768 ) );
  AOI22D0 U774 ( .A1(S_mag[20]), .A2(n700), .B1(n937), .B2(n699), .ZN(n651) );
  AOI22D0 U775 ( .A1(S_mag[22]), .A2(n701), .B1(S_mag[21]), .B2(n702), .ZN(
        n650) );
  CKND2D0 U776 ( .A1(n651), .A2(n650), .ZN(n652) );
  MUX2ND0 U777 ( .I0(n1029), .I1(n698), .S(n652), .ZN(
        \DP_OP_13J3_123_8774/n769 ) );
  AOI22D0 U778 ( .A1(n700), .A2(S_mag[19]), .B1(n699), .B2(n941), .ZN(n654) );
  AOI22D0 U779 ( .A1(S_mag[21]), .A2(n701), .B1(S_mag[20]), .B2(n702), .ZN(
        n653) );
  CKND2D0 U780 ( .A1(n654), .A2(n653), .ZN(n655) );
  MUX2ND0 U781 ( .I0(n1029), .I1(n698), .S(n655), .ZN(
        \DP_OP_13J3_123_8774/n770 ) );
  AOI22D0 U782 ( .A1(S_mag[18]), .A2(n700), .B1(n699), .B2(n945), .ZN(n657) );
  AOI22D0 U783 ( .A1(S_mag[20]), .A2(n701), .B1(n702), .B2(S_mag[19]), .ZN(
        n656) );
  CKND2D0 U784 ( .A1(n657), .A2(n656), .ZN(n658) );
  MUX2ND0 U785 ( .I0(n1029), .I1(n698), .S(n658), .ZN(
        \DP_OP_13J3_123_8774/n771 ) );
  AOI22D0 U786 ( .A1(S_mag[17]), .A2(n700), .B1(n699), .B2(n949), .ZN(n660) );
  AOI22D0 U787 ( .A1(S_mag[18]), .A2(n702), .B1(n701), .B2(S_mag[19]), .ZN(
        n659) );
  CKND2D0 U788 ( .A1(n660), .A2(n659), .ZN(n661) );
  MUX2ND0 U789 ( .I0(n1029), .I1(n698), .S(n661), .ZN(
        \DP_OP_13J3_123_8774/n772 ) );
  AOI22D0 U790 ( .A1(S_mag[16]), .A2(n700), .B1(n953), .B2(n699), .ZN(n663) );
  AOI22D0 U791 ( .A1(S_mag[17]), .A2(n702), .B1(S_mag[18]), .B2(n701), .ZN(
        n662) );
  CKND2D0 U792 ( .A1(n663), .A2(n662), .ZN(n664) );
  MUX2ND0 U793 ( .I0(n1029), .I1(n698), .S(n664), .ZN(
        \DP_OP_13J3_123_8774/n773 ) );
  AOI22D0 U794 ( .A1(S_mag[15]), .A2(n700), .B1(n957), .B2(n699), .ZN(n666) );
  AOI22D0 U795 ( .A1(S_mag[17]), .A2(n701), .B1(S_mag[16]), .B2(n702), .ZN(
        n665) );
  CKND2D0 U796 ( .A1(n666), .A2(n665), .ZN(n667) );
  MUX2ND0 U797 ( .I0(n1029), .I1(n698), .S(n667), .ZN(
        \DP_OP_13J3_123_8774/n774 ) );
  AOI22D0 U798 ( .A1(S_mag[14]), .A2(n700), .B1(n699), .B2(n961), .ZN(n669) );
  AOI22D0 U799 ( .A1(S_mag[15]), .A2(n702), .B1(S_mag[16]), .B2(n701), .ZN(
        n668) );
  CKND2D0 U800 ( .A1(n669), .A2(n668), .ZN(n670) );
  MUX2ND0 U801 ( .I0(n1029), .I1(n698), .S(n670), .ZN(
        \DP_OP_13J3_123_8774/n775 ) );
  AOI22D0 U802 ( .A1(S_mag[14]), .A2(n702), .B1(S_mag[15]), .B2(n701), .ZN(
        n671) );
  CKND2D0 U803 ( .A1(n672), .A2(n671), .ZN(n673) );
  MUX2ND0 U804 ( .I0(n1029), .I1(n698), .S(n673), .ZN(
        \DP_OP_13J3_123_8774/n776 ) );
  AOI22D0 U805 ( .A1(S_mag[12]), .A2(n700), .B1(n969), .B2(n699), .ZN(n675) );
  CKND2D0 U806 ( .A1(n675), .A2(n674), .ZN(n676) );
  MUX2ND0 U807 ( .I0(n1029), .I1(n698), .S(n676), .ZN(
        \DP_OP_13J3_123_8774/n777 ) );
  AOI22D0 U808 ( .A1(S_mag[13]), .A2(n701), .B1(n973), .B2(n699), .ZN(n678) );
  AOI22D0 U809 ( .A1(S_mag[12]), .A2(n702), .B1(S_mag[11]), .B2(n700), .ZN(
        n677) );
  CKND2D0 U810 ( .A1(n678), .A2(n677), .ZN(n679) );
  MUX2ND0 U811 ( .I0(n1029), .I1(n698), .S(n679), .ZN(
        \DP_OP_13J3_123_8774/n778 ) );
  AOI22D0 U812 ( .A1(S_mag[12]), .A2(n701), .B1(n977), .B2(n699), .ZN(n681) );
  AOI22D0 U813 ( .A1(S_mag[10]), .A2(n700), .B1(S_mag[11]), .B2(n702), .ZN(
        n680) );
  CKND2D0 U814 ( .A1(n681), .A2(n680), .ZN(n682) );
  MUX2ND0 U815 ( .I0(n1029), .I1(n698), .S(n682), .ZN(
        \DP_OP_13J3_123_8774/n779 ) );
  AOI22D0 U816 ( .A1(S_mag[9]), .A2(n700), .B1(n699), .B2(n981), .ZN(n684) );
  AOI22D0 U817 ( .A1(S_mag[10]), .A2(n702), .B1(S_mag[11]), .B2(n701), .ZN(
        n683) );
  MUX2ND0 U818 ( .I0(n1029), .I1(n698), .S(n685), .ZN(
        \DP_OP_13J3_123_8774/n780 ) );
  AOI22D0 U819 ( .A1(S_mag[8]), .A2(n700), .B1(n985), .B2(n699), .ZN(n687) );
  AOI22D0 U820 ( .A1(S_mag[9]), .A2(n702), .B1(S_mag[10]), .B2(n701), .ZN(n686) );
  CKND2D0 U821 ( .A1(n687), .A2(n686), .ZN(n688) );
  MUX2ND0 U822 ( .I0(n1029), .I1(n698), .S(n688), .ZN(
        \DP_OP_13J3_123_8774/n781 ) );
  AOI22D0 U823 ( .A1(S_mag[7]), .A2(n700), .B1(n989), .B2(n699), .ZN(n690) );
  AOI22D0 U824 ( .A1(S_mag[8]), .A2(n702), .B1(S_mag[9]), .B2(n701), .ZN(n689)
         );
  CKND2D0 U825 ( .A1(n690), .A2(n689), .ZN(n691) );
  MUX2ND0 U826 ( .I0(n1029), .I1(n698), .S(n691), .ZN(
        \DP_OP_13J3_123_8774/n782 ) );
  AOI22D0 U827 ( .A1(S_mag[6]), .A2(n700), .B1(n993), .B2(n699), .ZN(n693) );
  AOI22D0 U828 ( .A1(S_mag[7]), .A2(n702), .B1(S_mag[8]), .B2(n701), .ZN(n692)
         );
  CKND2D0 U829 ( .A1(n693), .A2(n692), .ZN(n694) );
  MUX2ND0 U830 ( .I0(n1029), .I1(n698), .S(n694), .ZN(
        \DP_OP_13J3_123_8774/n783 ) );
  AOI22D0 U831 ( .A1(S_mag[5]), .A2(n700), .B1(n997), .B2(n699), .ZN(n696) );
  AOI22D0 U832 ( .A1(S_mag[6]), .A2(n702), .B1(S_mag[7]), .B2(n701), .ZN(n695)
         );
  CKND2D0 U833 ( .A1(n696), .A2(n695), .ZN(n697) );
  MUX2ND0 U834 ( .I0(n1029), .I1(n698), .S(n697), .ZN(
        \DP_OP_13J3_123_8774/n784 ) );
  AOI22D0 U835 ( .A1(S_mag[4]), .A2(n700), .B1(n1002), .B2(n699), .ZN(n704) );
  AOI22D0 U836 ( .A1(S_mag[5]), .A2(n702), .B1(S_mag[6]), .B2(n701), .ZN(n703)
         );
  CKND2D0 U837 ( .A1(n704), .A2(n703), .ZN(n705) );
  MUX2ND0 U838 ( .I0(n1029), .I1(n698), .S(n705), .ZN(
        \DP_OP_13J3_123_8774/n785 ) );
  OAI22D0 U839 ( .A1(n933), .A2(n769), .B1(n928), .B2(n707), .ZN(n706) );
  MUX2ND0 U840 ( .I0(n709), .I1(n774), .S(n706), .ZN(
        \DP_OP_13J3_123_8774/n793 ) );
  OAI222D0 U841 ( .A1(n769), .A2(n930), .B1(n767), .B2(n933), .C1(n935), .C2(
        n707), .ZN(n708) );
  MUX2ND0 U842 ( .I0(n709), .I1(n774), .S(n708), .ZN(
        \DP_OP_13J3_123_8774/n794 ) );
  NR2D0 U843 ( .A1(n930), .A2(n767), .ZN(n711) );
  OAI22D0 U844 ( .A1(n933), .A2(n768), .B1(n846), .B2(n769), .ZN(n710) );
  MUX2ND0 U845 ( .I0(n774), .I1(n709), .S(n712), .ZN(
        \DP_OP_13J3_123_8774/n795 ) );
  NR2D0 U846 ( .A1(n846), .A2(n767), .ZN(n714) );
  AOI211D0 U847 ( .A1(n941), .A2(n772), .B(n714), .C(n713), .ZN(n715) );
  MUX2ND0 U848 ( .I0(n774), .I1(n709), .S(n715), .ZN(
        \DP_OP_13J3_123_8774/n796 ) );
  NR2D0 U849 ( .A1(n767), .A2(n850), .ZN(n717) );
  OAI22D0 U850 ( .A1(n846), .A2(n768), .B1(n854), .B2(n769), .ZN(n716) );
  AOI211D0 U851 ( .A1(n945), .A2(n772), .B(n717), .C(n716), .ZN(n718) );
  MUX2ND0 U852 ( .I0(n774), .I1(n709), .S(n718), .ZN(
        \DP_OP_13J3_123_8774/n797 ) );
  NR2D0 U853 ( .A1(n854), .A2(n767), .ZN(n720) );
  OAI22D0 U854 ( .A1(n858), .A2(n769), .B1(n768), .B2(n850), .ZN(n719) );
  AOI211D0 U855 ( .A1(n949), .A2(n772), .B(n720), .C(n719), .ZN(n721) );
  MUX2ND0 U856 ( .I0(n774), .I1(n709), .S(n721), .ZN(
        \DP_OP_13J3_123_8774/n798 ) );
  NR2D0 U857 ( .A1(n858), .A2(n767), .ZN(n723) );
  OAI22D0 U858 ( .A1(n862), .A2(n769), .B1(n854), .B2(n768), .ZN(n722) );
  AOI211D0 U859 ( .A1(n772), .A2(n953), .B(n723), .C(n722), .ZN(n724) );
  MUX2ND0 U860 ( .I0(n774), .I1(n709), .S(n724), .ZN(
        \DP_OP_13J3_123_8774/n799 ) );
  NR2D0 U861 ( .A1(n862), .A2(n767), .ZN(n726) );
  OAI22D0 U862 ( .A1(n866), .A2(n769), .B1(n858), .B2(n768), .ZN(n725) );
  AOI211D0 U863 ( .A1(n772), .A2(n957), .B(n726), .C(n725), .ZN(n727) );
  MUX2ND0 U864 ( .I0(n774), .I1(n709), .S(n727), .ZN(
        \DP_OP_13J3_123_8774/n800 ) );
  NR2D0 U865 ( .A1(n866), .A2(n767), .ZN(n729) );
  OAI22D0 U866 ( .A1(n870), .A2(n769), .B1(n862), .B2(n768), .ZN(n728) );
  AOI211D0 U867 ( .A1(n961), .A2(n772), .B(n729), .C(n728), .ZN(n730) );
  MUX2ND0 U868 ( .I0(n774), .I1(n709), .S(n730), .ZN(
        \DP_OP_13J3_123_8774/n801 ) );
  NR2D0 U869 ( .A1(n870), .A2(n767), .ZN(n732) );
  OAI22D0 U870 ( .A1(n874), .A2(n769), .B1(n866), .B2(n768), .ZN(n731) );
  AOI211D0 U871 ( .A1(n772), .A2(n965), .B(n732), .C(n731), .ZN(n733) );
  MUX2ND0 U872 ( .I0(n774), .I1(n709), .S(n733), .ZN(
        \DP_OP_13J3_123_8774/n802 ) );
  NR2D0 U873 ( .A1(n874), .A2(n767), .ZN(n735) );
  OAI22D0 U874 ( .A1(n870), .A2(n768), .B1(n878), .B2(n769), .ZN(n734) );
  AOI211D0 U875 ( .A1(n772), .A2(n969), .B(n735), .C(n734), .ZN(n736) );
  MUX2ND0 U876 ( .I0(n774), .I1(n709), .S(n736), .ZN(
        \DP_OP_13J3_123_8774/n803 ) );
  NR2D0 U877 ( .A1(n882), .A2(n769), .ZN(n738) );
  OAI22D0 U878 ( .A1(n874), .A2(n768), .B1(n878), .B2(n767), .ZN(n737) );
  AOI211D0 U879 ( .A1(n772), .A2(n973), .B(n738), .C(n737), .ZN(n739) );
  MUX2ND0 U880 ( .I0(n774), .I1(n709), .S(n739), .ZN(
        \DP_OP_13J3_123_8774/n804 ) );
  NR2D0 U881 ( .A1(n886), .A2(n769), .ZN(n741) );
  OAI22D0 U882 ( .A1(n878), .A2(n768), .B1(n882), .B2(n767), .ZN(n740) );
  AOI211D0 U883 ( .A1(n772), .A2(n977), .B(n741), .C(n740), .ZN(n742) );
  MUX2ND0 U884 ( .I0(n774), .I1(n709), .S(n742), .ZN(
        \DP_OP_13J3_123_8774/n805 ) );
  NR2D0 U885 ( .A1(n886), .A2(n767), .ZN(n744) );
  OAI22D0 U886 ( .A1(n890), .A2(n769), .B1(n882), .B2(n768), .ZN(n743) );
  MUX2ND0 U887 ( .I0(n774), .I1(n709), .S(n745), .ZN(
        \DP_OP_13J3_123_8774/n806 ) );
  NR2D0 U888 ( .A1(n890), .A2(n767), .ZN(n747) );
  OAI22D0 U889 ( .A1(n894), .A2(n769), .B1(n886), .B2(n768), .ZN(n746) );
  MUX2ND0 U890 ( .I0(n774), .I1(n709), .S(n748), .ZN(
        \DP_OP_13J3_123_8774/n807 ) );
  NR2D0 U891 ( .A1(n894), .A2(n767), .ZN(n750) );
  OAI22D0 U892 ( .A1(n898), .A2(n769), .B1(n890), .B2(n768), .ZN(n749) );
  AOI211D0 U893 ( .A1(n772), .A2(n989), .B(n750), .C(n749), .ZN(n751) );
  MUX2ND0 U894 ( .I0(n774), .I1(n709), .S(n751), .ZN(
        \DP_OP_13J3_123_8774/n808 ) );
  NR2D0 U895 ( .A1(n898), .A2(n767), .ZN(n753) );
  OAI22D0 U896 ( .A1(n902), .A2(n769), .B1(n894), .B2(n768), .ZN(n752) );
  AOI211D0 U897 ( .A1(n772), .A2(n993), .B(n753), .C(n752), .ZN(n754) );
  MUX2ND0 U898 ( .I0(n774), .I1(n709), .S(n754), .ZN(
        \DP_OP_13J3_123_8774/n809 ) );
  OAI22D0 U899 ( .A1(n906), .A2(n769), .B1(n898), .B2(n768), .ZN(n755) );
  AOI211D0 U900 ( .A1(n772), .A2(n997), .B(n756), .C(n755), .ZN(n757) );
  MUX2ND0 U901 ( .I0(n774), .I1(n709), .S(n757), .ZN(
        \DP_OP_13J3_123_8774/n810 ) );
  NR2D0 U902 ( .A1(n906), .A2(n767), .ZN(n759) );
  AOI211D0 U903 ( .A1(n772), .A2(n1002), .B(n759), .C(n758), .ZN(n760) );
  MUX2ND0 U904 ( .I0(n774), .I1(n709), .S(n760), .ZN(
        \DP_OP_13J3_123_8774/n811 ) );
  OAI22D0 U905 ( .A1(n919), .A2(n769), .B1(n906), .B2(n768), .ZN(n761) );
  AOI211D0 U906 ( .A1(n772), .A2(n909), .B(n762), .C(n761), .ZN(n763) );
  MUX2ND0 U907 ( .I0(n774), .I1(n709), .S(n763), .ZN(
        \DP_OP_13J3_123_8774/n812 ) );
  OAI22D0 U908 ( .A1(n917), .A2(n769), .B1(n911), .B2(n768), .ZN(n764) );
  AOI211D0 U909 ( .A1(n772), .A2(n914), .B(n765), .C(n764), .ZN(n766) );
  MUX2ND0 U910 ( .I0(n774), .I1(n709), .S(n766), .ZN(
        \DP_OP_13J3_123_8774/n813 ) );
  NR2D0 U911 ( .A1(n917), .A2(n767), .ZN(n771) );
  OAI22D0 U912 ( .A1(n921), .A2(n769), .B1(n919), .B2(n768), .ZN(n770) );
  AOI211D0 U913 ( .A1(n772), .A2(n924), .B(n771), .C(n770), .ZN(n773) );
  MUX2ND0 U914 ( .I0(n774), .I1(n709), .S(n773), .ZN(
        \DP_OP_13J3_123_8774/n814 ) );
  MUX2ND0 U915 ( .I0(n1030), .I1(n828), .S(n775), .ZN(
        \DP_OP_13J3_123_8774/n819 ) );
  INVD0 U916 ( .I(n832), .ZN(n777) );
  OAI222D0 U917 ( .A1(n778), .A2(n930), .B1(n777), .B2(n933), .C1(n935), .C2(
        n776), .ZN(n779) );
  MUX2ND0 U918 ( .I0(n1030), .I1(n828), .S(n779), .ZN(
        \DP_OP_13J3_123_8774/n820 ) );
  AOI22D0 U919 ( .A1(S_mag[20]), .A2(n830), .B1(n937), .B2(n829), .ZN(n781) );
  AOI22D0 U920 ( .A1(S_mag[22]), .A2(n831), .B1(S_mag[21]), .B2(n832), .ZN(
        n780) );
  CKND2D0 U921 ( .A1(n781), .A2(n780), .ZN(n782) );
  MUX2ND0 U922 ( .I0(n1030), .I1(n828), .S(n782), .ZN(
        \DP_OP_13J3_123_8774/n821 ) );
  AOI22D0 U923 ( .A1(n830), .A2(S_mag[19]), .B1(n829), .B2(n941), .ZN(n784) );
  AOI22D0 U924 ( .A1(S_mag[21]), .A2(n831), .B1(S_mag[20]), .B2(n832), .ZN(
        n783) );
  CKND2D0 U925 ( .A1(n784), .A2(n783), .ZN(n785) );
  MUX2ND0 U926 ( .I0(n1030), .I1(n828), .S(n785), .ZN(
        \DP_OP_13J3_123_8774/n822 ) );
  AOI22D0 U927 ( .A1(S_mag[18]), .A2(n830), .B1(n829), .B2(n945), .ZN(n787) );
  AOI22D0 U928 ( .A1(S_mag[20]), .A2(n831), .B1(n832), .B2(S_mag[19]), .ZN(
        n786) );
  CKND2D0 U929 ( .A1(n787), .A2(n786), .ZN(n788) );
  MUX2ND0 U930 ( .I0(n1030), .I1(n828), .S(n788), .ZN(
        \DP_OP_13J3_123_8774/n823 ) );
  AOI22D0 U931 ( .A1(S_mag[17]), .A2(n830), .B1(n829), .B2(n949), .ZN(n790) );
  AOI22D0 U932 ( .A1(S_mag[18]), .A2(n832), .B1(n831), .B2(S_mag[19]), .ZN(
        n789) );
  CKND2D0 U933 ( .A1(n790), .A2(n789), .ZN(n791) );
  MUX2ND0 U934 ( .I0(n1030), .I1(n828), .S(n791), .ZN(
        \DP_OP_13J3_123_8774/n824 ) );
  AOI22D0 U935 ( .A1(S_mag[16]), .A2(n830), .B1(n953), .B2(n829), .ZN(n793) );
  AOI22D0 U936 ( .A1(S_mag[17]), .A2(n832), .B1(S_mag[18]), .B2(n831), .ZN(
        n792) );
  MUX2ND0 U937 ( .I0(n1030), .I1(n828), .S(n794), .ZN(
        \DP_OP_13J3_123_8774/n825 ) );
  AOI22D0 U938 ( .A1(S_mag[15]), .A2(n830), .B1(n957), .B2(n829), .ZN(n796) );
  AOI22D0 U939 ( .A1(S_mag[17]), .A2(n831), .B1(S_mag[16]), .B2(n832), .ZN(
        n795) );
  CKND2D0 U940 ( .A1(n796), .A2(n795), .ZN(n797) );
  MUX2ND0 U941 ( .I0(n1030), .I1(n828), .S(n797), .ZN(
        \DP_OP_13J3_123_8774/n826 ) );
  AOI22D0 U942 ( .A1(S_mag[14]), .A2(n830), .B1(n829), .B2(n961), .ZN(n799) );
  AOI22D0 U943 ( .A1(S_mag[15]), .A2(n832), .B1(S_mag[16]), .B2(n831), .ZN(
        n798) );
  CKND2D0 U944 ( .A1(n799), .A2(n798), .ZN(n800) );
  MUX2ND0 U945 ( .I0(n1030), .I1(n828), .S(n800), .ZN(
        \DP_OP_13J3_123_8774/n827 ) );
  AOI22D0 U946 ( .A1(S_mag[13]), .A2(n830), .B1(n965), .B2(n829), .ZN(n802) );
  AOI22D0 U947 ( .A1(S_mag[14]), .A2(n832), .B1(S_mag[15]), .B2(n831), .ZN(
        n801) );
  CKND2D0 U948 ( .A1(n802), .A2(n801), .ZN(n803) );
  MUX2ND0 U949 ( .I0(n1030), .I1(n828), .S(n803), .ZN(
        \DP_OP_13J3_123_8774/n828 ) );
  AOI22D0 U950 ( .A1(S_mag[12]), .A2(n830), .B1(n969), .B2(n829), .ZN(n805) );
  AOI22D0 U951 ( .A1(S_mag[14]), .A2(n831), .B1(S_mag[13]), .B2(n832), .ZN(
        n804) );
  CKND2D0 U952 ( .A1(n805), .A2(n804), .ZN(n806) );
  MUX2ND0 U953 ( .I0(n1030), .I1(n828), .S(n806), .ZN(
        \DP_OP_13J3_123_8774/n829 ) );
  AOI22D0 U954 ( .A1(S_mag[13]), .A2(n831), .B1(n973), .B2(n829), .ZN(n808) );
  AOI22D0 U955 ( .A1(S_mag[12]), .A2(n832), .B1(S_mag[11]), .B2(n830), .ZN(
        n807) );
  CKND2D0 U956 ( .A1(n808), .A2(n807), .ZN(n809) );
  MUX2ND0 U957 ( .I0(n1030), .I1(n828), .S(n809), .ZN(
        \DP_OP_13J3_123_8774/n830 ) );
  AOI22D0 U958 ( .A1(S_mag[10]), .A2(n830), .B1(S_mag[11]), .B2(n832), .ZN(
        n810) );
  CKND2D0 U959 ( .A1(n811), .A2(n810), .ZN(n812) );
  MUX2ND0 U960 ( .I0(n1030), .I1(n828), .S(n812), .ZN(
        \DP_OP_13J3_123_8774/n831 ) );
  AOI22D0 U961 ( .A1(S_mag[9]), .A2(n830), .B1(n829), .B2(n981), .ZN(n814) );
  AOI22D0 U962 ( .A1(S_mag[10]), .A2(n832), .B1(S_mag[11]), .B2(n831), .ZN(
        n813) );
  CKND2D0 U963 ( .A1(n814), .A2(n813), .ZN(n815) );
  MUX2ND0 U964 ( .I0(n1030), .I1(n828), .S(n815), .ZN(
        \DP_OP_13J3_123_8774/n832 ) );
  AOI22D0 U965 ( .A1(S_mag[8]), .A2(n830), .B1(n985), .B2(n829), .ZN(n817) );
  AOI22D0 U966 ( .A1(S_mag[9]), .A2(n832), .B1(S_mag[10]), .B2(n831), .ZN(n816) );
  CKND2D0 U967 ( .A1(n817), .A2(n816), .ZN(n818) );
  MUX2ND0 U968 ( .I0(n1030), .I1(n828), .S(n818), .ZN(
        \DP_OP_13J3_123_8774/n833 ) );
  AOI22D0 U969 ( .A1(S_mag[7]), .A2(n830), .B1(n989), .B2(n829), .ZN(n820) );
  AOI22D0 U970 ( .A1(S_mag[8]), .A2(n832), .B1(S_mag[9]), .B2(n831), .ZN(n819)
         );
  CKND2D0 U971 ( .A1(n820), .A2(n819), .ZN(n821) );
  MUX2ND0 U972 ( .I0(n1030), .I1(n828), .S(n821), .ZN(
        \DP_OP_13J3_123_8774/n834 ) );
  AOI22D0 U973 ( .A1(S_mag[6]), .A2(n830), .B1(n993), .B2(n829), .ZN(n823) );
  AOI22D0 U974 ( .A1(S_mag[7]), .A2(n832), .B1(S_mag[8]), .B2(n831), .ZN(n822)
         );
  CKND2D0 U975 ( .A1(n823), .A2(n822), .ZN(n824) );
  MUX2ND0 U976 ( .I0(n1030), .I1(n828), .S(n824), .ZN(
        \DP_OP_13J3_123_8774/n835 ) );
  AOI22D0 U977 ( .A1(S_mag[5]), .A2(n830), .B1(n997), .B2(n829), .ZN(n826) );
  AOI22D0 U978 ( .A1(S_mag[6]), .A2(n832), .B1(S_mag[7]), .B2(n831), .ZN(n825)
         );
  CKND2D0 U979 ( .A1(n826), .A2(n825), .ZN(n827) );
  MUX2ND0 U980 ( .I0(n1030), .I1(n828), .S(n827), .ZN(
        \DP_OP_13J3_123_8774/n836 ) );
  AOI22D0 U981 ( .A1(S_mag[4]), .A2(n830), .B1(n1002), .B2(n829), .ZN(n834) );
  AOI22D0 U982 ( .A1(S_mag[5]), .A2(n832), .B1(S_mag[6]), .B2(n831), .ZN(n833)
         );
  CKND2D0 U983 ( .A1(n834), .A2(n833), .ZN(n835) );
  MUX2ND0 U984 ( .I0(n1030), .I1(n828), .S(n835), .ZN(
        \DP_OP_13J3_123_8774/n837 ) );
  OAI22D0 U985 ( .A1(n933), .A2(n920), .B1(n928), .B2(n837), .ZN(n836) );
  MUX2ND0 U986 ( .I0(n839), .I1(n927), .S(n836), .ZN(
        \DP_OP_13J3_123_8774/n845 ) );
  OAI222D0 U987 ( .A1(n920), .A2(n930), .B1(n916), .B2(n933), .C1(n935), .C2(
        n837), .ZN(n838) );
  MUX2ND0 U988 ( .I0(n839), .I1(n927), .S(n838), .ZN(
        \DP_OP_13J3_123_8774/n846 ) );
  NR2D0 U989 ( .A1(n930), .A2(n916), .ZN(n841) );
  OAI22D0 U990 ( .A1(n933), .A2(n918), .B1(n846), .B2(n920), .ZN(n840) );
  MUX2ND0 U991 ( .I0(n927), .I1(n839), .S(n842), .ZN(
        \DP_OP_13J3_123_8774/n847 ) );
  NR2D0 U992 ( .A1(n846), .A2(n916), .ZN(n844) );
  OAI22D0 U993 ( .A1(n930), .A2(n918), .B1(n920), .B2(n850), .ZN(n843) );
  AOI211D0 U994 ( .A1(n941), .A2(n925), .B(n844), .C(n843), .ZN(n845) );
  MUX2ND0 U995 ( .I0(n927), .I1(n839), .S(n845), .ZN(
        \DP_OP_13J3_123_8774/n848 ) );
  NR2D0 U996 ( .A1(n916), .A2(n850), .ZN(n848) );
  OAI22D0 U997 ( .A1(n846), .A2(n918), .B1(n854), .B2(n920), .ZN(n847) );
  AOI211D0 U998 ( .A1(n945), .A2(n925), .B(n848), .C(n847), .ZN(n849) );
  MUX2ND0 U999 ( .I0(n927), .I1(n839), .S(n849), .ZN(
        \DP_OP_13J3_123_8774/n849 ) );
  NR2D0 U1000 ( .A1(n854), .A2(n916), .ZN(n852) );
  OAI22D0 U1001 ( .A1(n858), .A2(n920), .B1(n918), .B2(n850), .ZN(n851) );
  AOI211D0 U1002 ( .A1(n949), .A2(n925), .B(n852), .C(n851), .ZN(n853) );
  MUX2ND0 U1003 ( .I0(n927), .I1(n839), .S(n853), .ZN(
        \DP_OP_13J3_123_8774/n850 ) );
  NR2D0 U1004 ( .A1(n858), .A2(n916), .ZN(n856) );
  OAI22D0 U1005 ( .A1(n862), .A2(n920), .B1(n854), .B2(n918), .ZN(n855) );
  AOI211D0 U1006 ( .A1(n925), .A2(n953), .B(n856), .C(n855), .ZN(n857) );
  MUX2ND0 U1007 ( .I0(n927), .I1(n839), .S(n857), .ZN(
        \DP_OP_13J3_123_8774/n851 ) );
  NR2D0 U1008 ( .A1(n862), .A2(n916), .ZN(n860) );
  OAI22D0 U1009 ( .A1(n866), .A2(n920), .B1(n858), .B2(n918), .ZN(n859) );
  AOI211D0 U1010 ( .A1(n925), .A2(n957), .B(n860), .C(n859), .ZN(n861) );
  MUX2ND0 U1011 ( .I0(n927), .I1(n839), .S(n861), .ZN(
        \DP_OP_13J3_123_8774/n852 ) );
  NR2D0 U1012 ( .A1(n866), .A2(n916), .ZN(n864) );
  OAI22D0 U1013 ( .A1(n870), .A2(n920), .B1(n862), .B2(n918), .ZN(n863) );
  AOI211D0 U1014 ( .A1(n961), .A2(n925), .B(n864), .C(n863), .ZN(n865) );
  MUX2ND0 U1015 ( .I0(n927), .I1(n839), .S(n865), .ZN(
        \DP_OP_13J3_123_8774/n853 ) );
  NR2D0 U1016 ( .A1(n870), .A2(n916), .ZN(n868) );
  OAI22D0 U1017 ( .A1(n874), .A2(n920), .B1(n866), .B2(n918), .ZN(n867) );
  AOI211D0 U1018 ( .A1(n925), .A2(n965), .B(n868), .C(n867), .ZN(n869) );
  MUX2ND0 U1019 ( .I0(n927), .I1(n839), .S(n869), .ZN(
        \DP_OP_13J3_123_8774/n854 ) );
  NR2D0 U1020 ( .A1(n874), .A2(n916), .ZN(n872) );
  OAI22D0 U1021 ( .A1(n870), .A2(n918), .B1(n878), .B2(n920), .ZN(n871) );
  AOI211D0 U1022 ( .A1(n925), .A2(n969), .B(n872), .C(n871), .ZN(n873) );
  MUX2ND0 U1023 ( .I0(n927), .I1(n839), .S(n873), .ZN(
        \DP_OP_13J3_123_8774/n855 ) );
  OAI22D0 U1024 ( .A1(n874), .A2(n918), .B1(n878), .B2(n916), .ZN(n875) );
  AOI211D0 U1025 ( .A1(n925), .A2(n973), .B(n876), .C(n875), .ZN(n877) );
  MUX2ND0 U1026 ( .I0(n927), .I1(n839), .S(n877), .ZN(
        \DP_OP_13J3_123_8774/n856 ) );
  NR2D0 U1027 ( .A1(n886), .A2(n920), .ZN(n880) );
  OAI22D0 U1028 ( .A1(n878), .A2(n918), .B1(n882), .B2(n916), .ZN(n879) );
  AOI211D0 U1029 ( .A1(n925), .A2(n977), .B(n880), .C(n879), .ZN(n881) );
  MUX2ND0 U1030 ( .I0(n927), .I1(n839), .S(n881), .ZN(
        \DP_OP_13J3_123_8774/n857 ) );
  OAI22D0 U1031 ( .A1(n890), .A2(n920), .B1(n882), .B2(n918), .ZN(n883) );
  AOI211D0 U1032 ( .A1(n981), .A2(n925), .B(n884), .C(n883), .ZN(n885) );
  MUX2ND0 U1033 ( .I0(n927), .I1(n839), .S(n885), .ZN(
        \DP_OP_13J3_123_8774/n858 ) );
  NR2D0 U1034 ( .A1(n890), .A2(n916), .ZN(n888) );
  OAI22D0 U1035 ( .A1(n894), .A2(n920), .B1(n886), .B2(n918), .ZN(n887) );
  AOI211D0 U1036 ( .A1(n925), .A2(n985), .B(n888), .C(n887), .ZN(n889) );
  MUX2ND0 U1037 ( .I0(n927), .I1(n839), .S(n889), .ZN(
        \DP_OP_13J3_123_8774/n859 ) );
  NR2D0 U1038 ( .A1(n894), .A2(n916), .ZN(n892) );
  OAI22D0 U1039 ( .A1(n898), .A2(n920), .B1(n890), .B2(n918), .ZN(n891) );
  AOI211D0 U1040 ( .A1(n925), .A2(n989), .B(n892), .C(n891), .ZN(n893) );
  MUX2ND0 U1041 ( .I0(n927), .I1(n839), .S(n893), .ZN(
        \DP_OP_13J3_123_8774/n860 ) );
  NR2D0 U1042 ( .A1(n898), .A2(n916), .ZN(n896) );
  OAI22D0 U1043 ( .A1(n902), .A2(n920), .B1(n894), .B2(n918), .ZN(n895) );
  MUX2ND0 U1044 ( .I0(n927), .I1(n839), .S(n897), .ZN(
        \DP_OP_13J3_123_8774/n861 ) );
  NR2D0 U1045 ( .A1(n902), .A2(n916), .ZN(n900) );
  OAI22D0 U1046 ( .A1(n906), .A2(n920), .B1(n898), .B2(n918), .ZN(n899) );
  AOI211D0 U1047 ( .A1(n925), .A2(n997), .B(n900), .C(n899), .ZN(n901) );
  MUX2ND0 U1048 ( .I0(n927), .I1(n839), .S(n901), .ZN(
        \DP_OP_13J3_123_8774/n862 ) );
  OAI22D0 U1049 ( .A1(n911), .A2(n920), .B1(n902), .B2(n918), .ZN(n903) );
  AOI211D0 U1050 ( .A1(n925), .A2(n1002), .B(n904), .C(n903), .ZN(n905) );
  MUX2ND0 U1051 ( .I0(n927), .I1(n839), .S(n905), .ZN(
        \DP_OP_13J3_123_8774/n863 ) );
  NR2D0 U1052 ( .A1(n911), .A2(n916), .ZN(n908) );
  OAI22D0 U1053 ( .A1(n919), .A2(n920), .B1(n906), .B2(n918), .ZN(n907) );
  AOI211D0 U1054 ( .A1(n925), .A2(n909), .B(n908), .C(n907), .ZN(n910) );
  MUX2ND0 U1055 ( .I0(n927), .I1(n839), .S(n910), .ZN(
        \DP_OP_13J3_123_8774/n864 ) );
  NR2D0 U1056 ( .A1(n919), .A2(n916), .ZN(n913) );
  OAI22D0 U1057 ( .A1(n917), .A2(n920), .B1(n911), .B2(n918), .ZN(n912) );
  AOI211D0 U1058 ( .A1(n925), .A2(n914), .B(n913), .C(n912), .ZN(n915) );
  MUX2ND0 U1059 ( .I0(n927), .I1(n839), .S(n915), .ZN(
        \DP_OP_13J3_123_8774/n865 ) );
  NR2D0 U1060 ( .A1(n917), .A2(n916), .ZN(n923) );
  OAI22D0 U1061 ( .A1(n921), .A2(n920), .B1(n919), .B2(n918), .ZN(n922) );
  AOI211D0 U1062 ( .A1(n925), .A2(n924), .B(n923), .C(n922), .ZN(n926) );
  MUX2ND0 U1063 ( .I0(n927), .I1(n839), .S(n926), .ZN(
        \DP_OP_13J3_123_8774/n866 ) );
  INVD0 U1064 ( .I(n1004), .ZN(n931) );
  OAI22D0 U1065 ( .A1(n931), .A2(n933), .B1(n934), .B2(n928), .ZN(n929) );
  MUX2ND0 U1066 ( .I0(n1028), .I1(n1001), .S(n929), .ZN(
        \DP_OP_13J3_123_8774/n871 ) );
  OAI222D0 U1067 ( .A1(n935), .A2(n934), .B1(n933), .B2(n932), .C1(n931), .C2(
        n930), .ZN(n936) );
  MUX2ND0 U1068 ( .I0(n1028), .I1(n1001), .S(n936), .ZN(
        \DP_OP_13J3_123_8774/n872 ) );
  AOI22D0 U1069 ( .A1(n1004), .A2(S_mag[20]), .B1(n1003), .B2(n937), .ZN(n939)
         );
  AOI22D0 U1070 ( .A1(n1006), .A2(S_mag[22]), .B1(n1005), .B2(S_mag[21]), .ZN(
        n938) );
  MUX2ND0 U1071 ( .I0(n1028), .I1(n1001), .S(n940), .ZN(
        \DP_OP_13J3_123_8774/n873 ) );
  AOI22D0 U1072 ( .A1(n1004), .A2(S_mag[19]), .B1(n1003), .B2(n941), .ZN(n943)
         );
  AOI22D0 U1073 ( .A1(n1006), .A2(S_mag[21]), .B1(n1005), .B2(S_mag[20]), .ZN(
        n942) );
  CKND2D0 U1074 ( .A1(n943), .A2(n942), .ZN(n944) );
  MUX2ND0 U1075 ( .I0(n1028), .I1(n1001), .S(n944), .ZN(
        \DP_OP_13J3_123_8774/n874 ) );
  AOI22D0 U1076 ( .A1(n1004), .A2(S_mag[18]), .B1(n1003), .B2(n945), .ZN(n947)
         );
  MUX2ND0 U1077 ( .I0(n1028), .I1(n1001), .S(n948), .ZN(
        \DP_OP_13J3_123_8774/n875 ) );
  AOI22D0 U1078 ( .A1(n1004), .A2(S_mag[17]), .B1(n1003), .B2(n949), .ZN(n951)
         );
  AOI22D0 U1079 ( .A1(n1006), .A2(S_mag[19]), .B1(n1005), .B2(S_mag[18]), .ZN(
        n950) );
  CKND2D0 U1080 ( .A1(n951), .A2(n950), .ZN(n952) );
  MUX2ND0 U1081 ( .I0(n1028), .I1(n1001), .S(n952), .ZN(
        \DP_OP_13J3_123_8774/n876 ) );
  AOI22D0 U1082 ( .A1(n1004), .A2(S_mag[16]), .B1(n1003), .B2(n953), .ZN(n955)
         );
  AOI22D0 U1083 ( .A1(n1006), .A2(S_mag[18]), .B1(n1005), .B2(S_mag[17]), .ZN(
        n954) );
  MUX2ND0 U1084 ( .I0(n1028), .I1(n1001), .S(n956), .ZN(
        \DP_OP_13J3_123_8774/n877 ) );
  AOI22D0 U1085 ( .A1(n1004), .A2(S_mag[15]), .B1(n1003), .B2(n957), .ZN(n959)
         );
  AOI22D0 U1086 ( .A1(n1006), .A2(S_mag[17]), .B1(n1005), .B2(S_mag[16]), .ZN(
        n958) );
  CKND2D0 U1087 ( .A1(n959), .A2(n958), .ZN(n960) );
  MUX2ND0 U1088 ( .I0(n1028), .I1(n1001), .S(n960), .ZN(
        \DP_OP_13J3_123_8774/n878 ) );
  AOI22D0 U1089 ( .A1(n1004), .A2(S_mag[14]), .B1(n1003), .B2(n961), .ZN(n963)
         );
  AOI22D0 U1090 ( .A1(n1006), .A2(S_mag[16]), .B1(n1005), .B2(S_mag[15]), .ZN(
        n962) );
  CKND2D0 U1091 ( .A1(n963), .A2(n962), .ZN(n964) );
  MUX2ND0 U1092 ( .I0(n1028), .I1(n1001), .S(n964), .ZN(
        \DP_OP_13J3_123_8774/n879 ) );
  AOI22D0 U1093 ( .A1(n1004), .A2(S_mag[13]), .B1(n1003), .B2(n965), .ZN(n967)
         );
  AOI22D0 U1094 ( .A1(n1006), .A2(S_mag[15]), .B1(n1005), .B2(S_mag[14]), .ZN(
        n966) );
  CKND2D0 U1095 ( .A1(n967), .A2(n966), .ZN(n968) );
  MUX2ND0 U1096 ( .I0(n1028), .I1(n1001), .S(n968), .ZN(
        \DP_OP_13J3_123_8774/n880 ) );
  AOI22D0 U1097 ( .A1(n1004), .A2(S_mag[12]), .B1(n1003), .B2(n969), .ZN(n971)
         );
  AOI22D0 U1098 ( .A1(n1006), .A2(S_mag[14]), .B1(n1005), .B2(S_mag[13]), .ZN(
        n970) );
  CKND2D0 U1099 ( .A1(n971), .A2(n970), .ZN(n972) );
  MUX2ND0 U1100 ( .I0(n1028), .I1(n1001), .S(n972), .ZN(
        \DP_OP_13J3_123_8774/n881 ) );
  AOI22D0 U1101 ( .A1(n1006), .A2(S_mag[13]), .B1(n1003), .B2(n973), .ZN(n975)
         );
  AOI22D0 U1102 ( .A1(n1005), .A2(S_mag[12]), .B1(n1004), .B2(S_mag[11]), .ZN(
        n974) );
  CKND2D0 U1103 ( .A1(n975), .A2(n974), .ZN(n976) );
  MUX2ND0 U1104 ( .I0(n1028), .I1(n1001), .S(n976), .ZN(
        \DP_OP_13J3_123_8774/n882 ) );
  AOI22D0 U1105 ( .A1(n1006), .A2(S_mag[12]), .B1(n1003), .B2(n977), .ZN(n979)
         );
  AOI22D0 U1106 ( .A1(n1005), .A2(S_mag[11]), .B1(n1004), .B2(S_mag[10]), .ZN(
        n978) );
  CKND2D0 U1107 ( .A1(n979), .A2(n978), .ZN(n980) );
  MUX2ND0 U1108 ( .I0(n1028), .I1(n1001), .S(n980), .ZN(
        \DP_OP_13J3_123_8774/n883 ) );
  AOI22D0 U1109 ( .A1(n1004), .A2(S_mag[9]), .B1(n1003), .B2(n981), .ZN(n983)
         );
  AOI22D0 U1110 ( .A1(n1006), .A2(S_mag[11]), .B1(n1005), .B2(S_mag[10]), .ZN(
        n982) );
  CKND2D0 U1111 ( .A1(n983), .A2(n982), .ZN(n984) );
  MUX2ND0 U1112 ( .I0(n1028), .I1(n1001), .S(n984), .ZN(
        \DP_OP_13J3_123_8774/n884 ) );
  AOI22D0 U1113 ( .A1(n1004), .A2(S_mag[8]), .B1(n1003), .B2(n985), .ZN(n987)
         );
  AOI22D0 U1114 ( .A1(n1006), .A2(S_mag[10]), .B1(n1005), .B2(S_mag[9]), .ZN(
        n986) );
  CKND2D0 U1115 ( .A1(n987), .A2(n986), .ZN(n988) );
  MUX2ND0 U1116 ( .I0(n1028), .I1(n1001), .S(n988), .ZN(
        \DP_OP_13J3_123_8774/n885 ) );
  AOI22D0 U1117 ( .A1(n1004), .A2(S_mag[7]), .B1(n1003), .B2(n989), .ZN(n991)
         );
  AOI22D0 U1118 ( .A1(n1006), .A2(S_mag[9]), .B1(n1005), .B2(S_mag[8]), .ZN(
        n990) );
  CKND2D0 U1119 ( .A1(n991), .A2(n990), .ZN(n992) );
  MUX2ND0 U1120 ( .I0(n1028), .I1(n1001), .S(n992), .ZN(
        \DP_OP_13J3_123_8774/n886 ) );
  AOI22D0 U1121 ( .A1(n1004), .A2(S_mag[6]), .B1(n1003), .B2(n993), .ZN(n995)
         );
  CKND2D0 U1122 ( .A1(n995), .A2(n994), .ZN(n996) );
  MUX2ND0 U1123 ( .I0(n1028), .I1(n1001), .S(n996), .ZN(
        \DP_OP_13J3_123_8774/n887 ) );
  AOI22D0 U1124 ( .A1(n1004), .A2(S_mag[5]), .B1(n1003), .B2(n997), .ZN(n999)
         );
  AOI22D0 U1125 ( .A1(n1006), .A2(S_mag[7]), .B1(n1005), .B2(S_mag[6]), .ZN(
        n998) );
  CKND2D0 U1126 ( .A1(n999), .A2(n998), .ZN(n1000) );
  MUX2ND0 U1127 ( .I0(n1028), .I1(n1001), .S(n1000), .ZN(
        \DP_OP_13J3_123_8774/n888 ) );
  AOI22D0 U1128 ( .A1(n1004), .A2(S_mag[4]), .B1(n1003), .B2(n1002), .ZN(n1008) );
  AOI22D0 U1129 ( .A1(n1006), .A2(S_mag[6]), .B1(n1005), .B2(S_mag[5]), .ZN(
        n1007) );
  MUX2ND0 U1130 ( .I0(n1028), .I1(n1001), .S(n1009), .ZN(
        \DP_OP_13J3_123_8774/n889 ) );
  AOI22D0 U1131 ( .A1(bit_pos[0]), .A2(n72), .B1(n1011), .B2(n1010), .ZN(n74)
         );
  INR2D0 U1132 ( .A1(n1012), .B1(n1016), .ZN(n1021) );
  AO22D0 U1133 ( .A1(n1027), .A2(n1021), .B1(Q_mag[22]), .B2(n1025), .Z(n68)
         );
  INR2D0 U1134 ( .A1(n1013), .B1(n1016), .ZN(n1026) );
  AO22D0 U1135 ( .A1(n1015), .A2(n1026), .B1(Q_mag[1]), .B2(n1025), .Z(n66) );
  AO22D0 U1136 ( .A1(Q_mag[2]), .A2(n1025), .B1(n1015), .B2(n1021), .Z(n65) );
  NR2D0 U1137 ( .A1(n1014), .A2(n1016), .ZN(n1022) );
  AO22D0 U1138 ( .A1(n1015), .A2(n1022), .B1(Q_mag[3]), .B2(n1025), .Z(n64) );
  INR2D0 U1139 ( .A1(n1017), .B1(n1016), .ZN(n1024) );
  AO22D0 U1140 ( .A1(n1018), .A2(n1024), .B1(Q_mag[4]), .B2(n1025), .Z(n63) );
  AO22D0 U1141 ( .A1(Q_mag[5]), .A2(n1025), .B1(n1018), .B2(n1026), .Z(n62) );
  AO22D0 U1142 ( .A1(n1018), .A2(n1021), .B1(Q_mag[6]), .B2(n1025), .Z(n61) );
  AO22D0 U1143 ( .A1(n1018), .A2(n1022), .B1(Q_mag[7]), .B2(n1025), .Z(n60) );
  AO22D0 U1144 ( .A1(n1019), .A2(n1024), .B1(Q_mag[8]), .B2(n1025), .Z(n59) );
  AO22D0 U1145 ( .A1(n1019), .A2(n1026), .B1(Q_mag[9]), .B2(n1025), .Z(n58) );
  AO22D0 U1146 ( .A1(n1021), .A2(n1019), .B1(Q_mag[10]), .B2(n1025), .Z(n57)
         );
  AO22D0 U1147 ( .A1(n1019), .A2(n1022), .B1(Q_mag[11]), .B2(n1025), .Z(n56)
         );
  AO22D0 U1148 ( .A1(n1020), .A2(n1024), .B1(Q_mag[12]), .B2(n1025), .Z(n55)
         );
  AO22D0 U1149 ( .A1(n1020), .A2(n1026), .B1(Q_mag[13]), .B2(n1025), .Z(n54)
         );
  AO22D0 U1150 ( .A1(n1021), .A2(n1020), .B1(Q_mag[14]), .B2(n1025), .Z(n53)
         );
  AO22D0 U1151 ( .A1(n1020), .A2(n1022), .B1(Q_mag[15]), .B2(n1025), .Z(n52)
         );
  AO22D0 U1152 ( .A1(n1023), .A2(n1024), .B1(Q_mag[16]), .B2(n1025), .Z(n51)
         );
  AO22D0 U1153 ( .A1(n1023), .A2(n1026), .B1(Q_mag[17]), .B2(n1025), .Z(n50)
         );
  AO22D0 U1154 ( .A1(n1021), .A2(n1023), .B1(Q_mag[18]), .B2(n1025), .Z(n49)
         );
  AO22D0 U1155 ( .A1(n1023), .A2(n1022), .B1(Q_mag[19]), .B2(n1025), .Z(n48)
         );
  AO22D0 U1156 ( .A1(n1027), .A2(n1024), .B1(Q_mag[20]), .B2(n1025), .Z(n47)
         );
  AO22D0 U1157 ( .A1(n1027), .A2(n1026), .B1(Q_mag[21]), .B2(n1025), .Z(n46)
         );
  CMPE42D1 U1158 ( .A(\DP_OP_13J3_123_8774/n445 ), .B(
        \DP_OP_13J3_123_8774/n439 ), .C(\DP_OP_13J3_123_8774/n797 ), .CIX(
        \DP_OP_13J3_123_8774/n820 ), .D(\DP_OP_13J3_123_8774/n441 ), .CO(
        \DP_OP_13J3_123_8774/n435 ), .COX(\DP_OP_13J3_123_8774/n434 ), .S(
        \DP_OP_13J3_123_8774/n436 ) );
  CMPE42D1 U1159 ( .A(\DP_OP_13J3_123_8774/n507 ), .B(
        \DP_OP_13J3_123_8774/n499 ), .C(\DP_OP_13J3_123_8774/n850 ), .CIX(
        \DP_OP_13J3_123_8774/n873 ), .D(\DP_OP_13J3_123_8774/n503 ), .CO(
        \DP_OP_13J3_123_8774/n495 ), .COX(\DP_OP_13J3_123_8774/n494 ), .S(
        \DP_OP_13J3_123_8774/n496 ) );
  CMPE42D1 U1160 ( .A(\DP_OP_13J3_123_8774/n472 ), .B(
        \DP_OP_13J3_123_8774/n464 ), .C(\DP_OP_13J3_123_8774/n823 ), .CIX(
        \DP_OP_13J3_123_8774/n846 ), .D(\DP_OP_13J3_123_8774/n468 ), .CO(
        \DP_OP_13J3_123_8774/n460 ), .COX(\DP_OP_13J3_123_8774/n459 ), .S(
        \DP_OP_13J3_123_8774/n461 ) );
  CMPE42D1 U1161 ( .A(\DP_OP_13J3_123_8774/n448 ), .B(
        \DP_OP_13J3_123_8774/n455 ), .C(\DP_OP_13J3_123_8774/n752 ), .CIX(
        \DP_OP_13J3_123_8774/n775 ), .D(\DP_OP_13J3_123_8774/n452 ), .CO(
        \DP_OP_13J3_123_8774/n445 ), .COX(\DP_OP_13J3_123_8774/n444 ), .S(
        \DP_OP_13J3_123_8774/n446 ) );
  CMPE42D1 U1162 ( .A(\DP_OP_13J3_123_8774/n475 ), .B(
        \DP_OP_13J3_123_8774/n483 ), .C(\DP_OP_13J3_123_8774/n778 ), .CIX(
        \DP_OP_13J3_123_8774/n801 ), .D(\DP_OP_13J3_123_8774/n479 ), .CO(
        \DP_OP_13J3_123_8774/n472 ), .COX(\DP_OP_13J3_123_8774/n471 ), .S(
        \DP_OP_13J3_123_8774/n473 ) );
  CMPE42D1 U1163 ( .A(n1030), .B(\DP_OP_13J3_123_8774/n432 ), .C(
        \DP_OP_13J3_123_8774/n727 ), .CIX(\DP_OP_13J3_123_8774/n749 ), .D(
        \DP_OP_13J3_123_8774/n429 ), .CO(\DP_OP_13J3_123_8774/n424 ), .COX(
        \DP_OP_13J3_123_8774/n413 ), .S(\DP_OP_13J3_123_8774/n425 ) );
  CMPE42D1 U1164 ( .A(n1028), .B(n1032), .C(\DP_OP_13J3_123_8774/n732 ), .CIX(
        \DP_OP_13J3_123_8774/n755 ), .D(\DP_OP_13J3_123_8774/n482 ), .CO(
        \DP_OP_13J3_123_8774/n474 ), .COX(\DP_OP_13J3_123_8774/n457 ), .S(
        \DP_OP_13J3_123_8774/n475 ) );
  CMPE42D1 U1165 ( .A(\DP_OP_13J3_123_8774/n736 ), .B(
        \DP_OP_13J3_123_8774/n759 ), .C(\DP_OP_13J3_123_8774/n518 ), .CIX(
        \DP_OP_13J3_123_8774/n519 ), .D(\DP_OP_13J3_123_8774/n782 ), .CO(
        \DP_OP_13J3_123_8774/n510 ), .COX(\DP_OP_13J3_123_8774/n509 ), .S(
        \DP_OP_13J3_123_8774/n511 ) );
  CMPE42D1 U1166 ( .A(\DP_OP_13J3_123_8774/n511 ), .B(
        \DP_OP_13J3_123_8774/n805 ), .C(\DP_OP_13J3_123_8774/n515 ), .CIX(
        \DP_OP_13J3_123_8774/n516 ), .D(\DP_OP_13J3_123_8774/n828 ), .CO(
        \DP_OP_13J3_123_8774/n507 ), .COX(\DP_OP_13J3_123_8774/n506 ), .S(
        \DP_OP_13J3_123_8774/n508 ) );
  CMPE42D1 U1167 ( .A(\DP_OP_13J3_123_8774/n723 ), .B(
        \DP_OP_13J3_123_8774/n403 ), .C(\DP_OP_13J3_123_8774/n745 ), .CIX(
        \DP_OP_13J3_123_8774/n768 ), .D(\DP_OP_13J3_123_8774/n404 ), .CO(
        \DP_OP_13J3_123_8774/n401 ), .COX(\DP_OP_13J3_123_8774/n400 ), .S(
        \DP_OP_13J3_123_8774/n402 ) );
  CMPE42D1 U1168 ( .A(\DP_OP_13J3_123_8774/n424 ), .B(
        \DP_OP_13J3_123_8774/n419 ), .C(\DP_OP_13J3_123_8774/n771 ), .CIX(
        \DP_OP_13J3_123_8774/n794 ), .D(\DP_OP_13J3_123_8774/n421 ), .CO(
        \DP_OP_13J3_123_8774/n416 ), .COX(\DP_OP_13J3_123_8774/n415 ), .S(
        \DP_OP_13J3_123_8774/n417 ) );
  CMPE42D1 U1169 ( .A(\DP_OP_13J3_123_8774/n446 ), .B(
        \DP_OP_13J3_123_8774/n453 ), .C(\DP_OP_13J3_123_8774/n798 ), .CIX(
        \DP_OP_13J3_123_8774/n821 ), .D(\DP_OP_13J3_123_8774/n449 ), .CO(
        \DP_OP_13J3_123_8774/n442 ), .COX(\DP_OP_13J3_123_8774/n441 ), .S(
        \DP_OP_13J3_123_8774/n443 ) );
  CMPE42D1 U1170 ( .A(\DP_OP_13J3_123_8774/n773 ), .B(
        \DP_OP_13J3_123_8774/n431 ), .C(\DP_OP_13J3_123_8774/n434 ), .CIX(
        \DP_OP_13J3_123_8774/n819 ), .D(\DP_OP_13J3_123_8774/n796 ), .CO(
        \DP_OP_13J3_123_8774/n427 ), .COX(\DP_OP_13J3_123_8774/n426 ), .S(
        \DP_OP_13J3_123_8774/n428 ) );
  CMPE42D1 U1171 ( .A(\DP_OP_13J3_123_8774/n403 ), .B(
        \DP_OP_13J3_123_8774/n722 ), .C(\DP_OP_13J3_123_8774/n400 ), .CIX(
        \DP_OP_13J3_123_8774/n767 ), .D(\DP_OP_13J3_123_8774/n744 ), .CO(
        \DP_OP_13J3_123_8774/n396 ), .COX(\DP_OP_13J3_123_8774/n395 ), .S(
        \DP_OP_13J3_123_8774/n397 ) );
  CMPE42D1 U1172 ( .A(\DP_OP_13J3_123_8774/n473 ), .B(
        \DP_OP_13J3_123_8774/n480 ), .C(\DP_OP_13J3_123_8774/n824 ), .CIX(
        \DP_OP_13J3_123_8774/n847 ), .D(\DP_OP_13J3_123_8774/n476 ), .CO(
        \DP_OP_13J3_123_8774/n469 ), .COX(\DP_OP_13J3_123_8774/n468 ), .S(
        \DP_OP_13J3_123_8774/n470 ) );
  CMPE42D1 U1173 ( .A(\DP_OP_13J3_123_8774/n425 ), .B(
        \DP_OP_13J3_123_8774/n430 ), .C(\DP_OP_13J3_123_8774/n772 ), .CIX(
        \DP_OP_13J3_123_8774/n795 ), .D(\DP_OP_13J3_123_8774/n426 ), .CO(
        \DP_OP_13J3_123_8774/n422 ), .COX(\DP_OP_13J3_123_8774/n421 ), .S(
        \DP_OP_13J3_123_8774/n423 ) );
  CMPE42D1 U1174 ( .A(\DP_OP_13J3_123_8774/n799 ), .B(
        \DP_OP_13J3_123_8774/n454 ), .C(\DP_OP_13J3_123_8774/n459 ), .CIX(
        \DP_OP_13J3_123_8774/n845 ), .D(\DP_OP_13J3_123_8774/n822 ), .CO(
        \DP_OP_13J3_123_8774/n450 ), .COX(\DP_OP_13J3_123_8774/n449 ), .S(
        \DP_OP_13J3_123_8774/n451 ) );
  CMPE42D1 U1175 ( .A(n1031), .B(\DP_OP_13J3_123_8774/n733 ), .C(
        \DP_OP_13J3_123_8774/n491 ), .CIX(\DP_OP_13J3_123_8774/n492 ), .D(
        \DP_OP_13J3_123_8774/n756 ), .CO(\DP_OP_13J3_123_8774/n483 ), .COX(
        \DP_OP_13J3_123_8774/n482 ), .S(\DP_OP_13J3_123_8774/n484 ) );
  CMPE42D1 U1176 ( .A(\DP_OP_13J3_123_8774/n779 ), .B(
        \DP_OP_13J3_123_8774/n484 ), .C(\DP_OP_13J3_123_8774/n488 ), .CIX(
        \DP_OP_13J3_123_8774/n489 ), .D(\DP_OP_13J3_123_8774/n802 ), .CO(
        \DP_OP_13J3_123_8774/n480 ), .COX(\DP_OP_13J3_123_8774/n479 ), .S(
        \DP_OP_13J3_123_8774/n481 ) );
  CMPE42D1 U1177 ( .A(\DP_OP_13J3_123_8774/n465 ), .B(
        \DP_OP_13J3_123_8774/n456 ), .C(\DP_OP_13J3_123_8774/n462 ), .CIX(
        \DP_OP_13J3_123_8774/n463 ), .D(\DP_OP_13J3_123_8774/n776 ), .CO(
        \DP_OP_13J3_123_8774/n453 ), .COX(\DP_OP_13J3_123_8774/n452 ), .S(
        \DP_OP_13J3_123_8774/n454 ) );
  CMPE42D1 U1178 ( .A(\DP_OP_13J3_123_8774/n440 ), .B(
        \DP_OP_13J3_123_8774/n728 ), .C(\DP_OP_13J3_123_8774/n437 ), .CIX(
        \DP_OP_13J3_123_8774/n438 ), .D(\DP_OP_13J3_123_8774/n750 ), .CO(
        \DP_OP_13J3_123_8774/n430 ), .COX(\DP_OP_13J3_123_8774/n429 ), .S(
        \DP_OP_13J3_123_8774/n431 ) );
  CMPE42D1 U1179 ( .A(\DP_OP_13J3_123_8774/n826 ), .B(
        \DP_OP_13J3_123_8774/n490 ), .C(\DP_OP_13J3_123_8774/n494 ), .CIX(
        \DP_OP_13J3_123_8774/n872 ), .D(\DP_OP_13J3_123_8774/n849 ), .CO(
        \DP_OP_13J3_123_8774/n486 ), .COX(\DP_OP_13J3_123_8774/n485 ), .S(
        \DP_OP_13J3_123_8774/n487 ) );
  CMPE42D1 U1180 ( .A(n1029), .B(\DP_OP_13J3_123_8774/n398 ), .C(
        \DP_OP_13J3_123_8774/n721 ), .CIX(\DP_OP_13J3_123_8774/n743 ), .D(
        \DP_OP_13J3_123_8774/n395 ), .CO(\DP_OP_13J3_123_8774/n393 ), .COX(
        \DP_OP_13J3_123_8774/n388 ), .S(\DP_OP_13J3_123_8774/n394 ) );
  CMPE42D1 U1181 ( .A(\DP_OP_13J3_123_8774/n747 ), .B(
        \DP_OP_13J3_123_8774/n412 ), .C(\DP_OP_13J3_123_8774/n415 ), .CIX(
        \DP_OP_13J3_123_8774/n793 ), .D(\DP_OP_13J3_123_8774/n770 ), .CO(
        \DP_OP_13J3_123_8774/n409 ), .COX(\DP_OP_13J3_123_8774/n408 ), .S(
        \DP_OP_13J3_123_8774/n410 ) );
  CMPE42D1 U1182 ( .A(\DP_OP_13J3_123_8774/n825 ), .B(
        \DP_OP_13J3_123_8774/n481 ), .C(\DP_OP_13J3_123_8774/n485 ), .CIX(
        \DP_OP_13J3_123_8774/n871 ), .D(\DP_OP_13J3_123_8774/n848 ), .CO(
        \DP_OP_13J3_123_8774/n477 ), .COX(\DP_OP_13J3_123_8774/n476 ), .S(
        \DP_OP_13J3_123_8774/n478 ) );
  CMPE42D1 U1183 ( .A(n1031), .B(\DP_OP_13J3_123_8774/n735 ), .C(
        \DP_OP_13J3_123_8774/n758 ), .CIX(\DP_OP_13J3_123_8774/n781 ), .D(
        \DP_OP_13J3_123_8774/n509 ), .CO(\DP_OP_13J3_123_8774/n501 ), .COX(
        \DP_OP_13J3_123_8774/n500 ), .S(\DP_OP_13J3_123_8774/n502 ) );
  CMPE42D1 U1184 ( .A(\DP_OP_13J3_123_8774/n510 ), .B(
        \DP_OP_13J3_123_8774/n502 ), .C(\DP_OP_13J3_123_8774/n804 ), .CIX(
        \DP_OP_13J3_123_8774/n827 ), .D(\DP_OP_13J3_123_8774/n506 ), .CO(
        \DP_OP_13J3_123_8774/n498 ), .COX(\DP_OP_13J3_123_8774/n497 ), .S(
        \DP_OP_13J3_123_8774/n499 ) );
  CMPE42D1 U1185 ( .A(\DP_OP_13J3_123_8774/n447 ), .B(
        \DP_OP_13J3_123_8774/n440 ), .C(\DP_OP_13J3_123_8774/n751 ), .CIX(
        \DP_OP_13J3_123_8774/n774 ), .D(\DP_OP_13J3_123_8774/n444 ), .CO(
        \DP_OP_13J3_123_8774/n438 ), .COX(\DP_OP_13J3_123_8774/n437 ), .S(
        \DP_OP_13J3_123_8774/n439 ) );
  CMPE42D1 U1186 ( .A(\DP_OP_13J3_123_8774/n474 ), .B(
        \DP_OP_13J3_123_8774/n466 ), .C(\DP_OP_13J3_123_8774/n777 ), .CIX(
        \DP_OP_13J3_123_8774/n800 ), .D(\DP_OP_13J3_123_8774/n471 ), .CO(
        \DP_OP_13J3_123_8774/n463 ), .COX(\DP_OP_13J3_123_8774/n462 ), .S(
        \DP_OP_13J3_123_8774/n464 ) );
  CMPE42D1 U1187 ( .A(\DP_OP_13J3_123_8774/n584 ), .B(
        \DP_OP_13J3_123_8774/n813 ), .C(\DP_OP_13J3_123_8774/n588 ), .CIX(
        \DP_OP_13J3_123_8774/n589 ), .D(\DP_OP_13J3_123_8774/n836 ), .CO(
        \DP_OP_13J3_123_8774/n581 ), .COX(\DP_OP_13J3_123_8774/n580 ), .S(
        \DP_OP_13J3_123_8774/n582 ) );
  CMPE42D1 U1188 ( .A(\DP_OP_13J3_123_8774/n576 ), .B(
        \DP_OP_13J3_123_8774/n812 ), .C(\DP_OP_13J3_123_8774/n580 ), .CIX(
        \DP_OP_13J3_123_8774/n581 ), .D(\DP_OP_13J3_123_8774/n835 ), .CO(
        \DP_OP_13J3_123_8774/n573 ), .COX(\DP_OP_13J3_123_8774/n572 ), .S(
        \DP_OP_13J3_123_8774/n574 ) );
  CMPE42D1 U1189 ( .A(\DP_OP_13J3_123_8774/n566 ), .B(
        \DP_OP_13J3_123_8774/n811 ), .C(\DP_OP_13J3_123_8774/n572 ), .CIX(
        \DP_OP_13J3_123_8774/n573 ), .D(\DP_OP_13J3_123_8774/n834 ), .CO(
        \DP_OP_13J3_123_8774/n563 ), .COX(\DP_OP_13J3_123_8774/n562 ), .S(
        \DP_OP_13J3_123_8774/n564 ) );
  CMPE42D1 U1190 ( .A(\DP_OP_13J3_123_8774/n738 ), .B(
        \DP_OP_13J3_123_8774/n761 ), .C(\DP_OP_13J3_123_8774/n536 ), .CIX(
        \DP_OP_13J3_123_8774/n537 ), .D(\DP_OP_13J3_123_8774/n784 ), .CO(
        \DP_OP_13J3_123_8774/n528 ), .COX(\DP_OP_13J3_123_8774/n527 ), .S(
        \DP_OP_13J3_123_8774/n529 ) );
  CMPE42D1 U1191 ( .A(\DP_OP_13J3_123_8774/n556 ), .B(
        \DP_OP_13J3_123_8774/n810 ), .C(\DP_OP_13J3_123_8774/n562 ), .CIX(
        \DP_OP_13J3_123_8774/n563 ), .D(\DP_OP_13J3_123_8774/n833 ), .CO(
        \DP_OP_13J3_123_8774/n553 ), .COX(\DP_OP_13J3_123_8774/n552 ), .S(
        \DP_OP_13J3_123_8774/n554 ) );
  CMPE42D1 U1192 ( .A(\DP_OP_13J3_123_8774/n737 ), .B(
        \DP_OP_13J3_123_8774/n760 ), .C(\DP_OP_13J3_123_8774/n527 ), .CIX(
        \DP_OP_13J3_123_8774/n528 ), .D(\DP_OP_13J3_123_8774/n783 ), .CO(
        \DP_OP_13J3_123_8774/n519 ), .COX(\DP_OP_13J3_123_8774/n518 ), .S(
        \DP_OP_13J3_123_8774/n520 ) );
  CMPE42D1 U1193 ( .A(\DP_OP_13J3_123_8774/n546 ), .B(
        \DP_OP_13J3_123_8774/n809 ), .C(\DP_OP_13J3_123_8774/n552 ), .CIX(
        \DP_OP_13J3_123_8774/n553 ), .D(\DP_OP_13J3_123_8774/n832 ), .CO(
        \DP_OP_13J3_123_8774/n543 ), .COX(\DP_OP_13J3_123_8774/n542 ), .S(
        \DP_OP_13J3_123_8774/n544 ) );
  CMPE42D1 U1194 ( .A(\DP_OP_13J3_123_8774/n538 ), .B(
        \DP_OP_13J3_123_8774/n808 ), .C(\DP_OP_13J3_123_8774/n542 ), .CIX(
        \DP_OP_13J3_123_8774/n543 ), .D(\DP_OP_13J3_123_8774/n831 ), .CO(
        \DP_OP_13J3_123_8774/n534 ), .COX(\DP_OP_13J3_123_8774/n533 ), .S(
        \DP_OP_13J3_123_8774/n535 ) );
  CMPE42D1 U1195 ( .A(\DP_OP_13J3_123_8774/n529 ), .B(
        \DP_OP_13J3_123_8774/n807 ), .C(\DP_OP_13J3_123_8774/n533 ), .CIX(
        \DP_OP_13J3_123_8774/n534 ), .D(\DP_OP_13J3_123_8774/n830 ), .CO(
        \DP_OP_13J3_123_8774/n525 ), .COX(\DP_OP_13J3_123_8774/n524 ), .S(
        \DP_OP_13J3_123_8774/n526 ) );
  CMPE42D1 U1196 ( .A(n1031), .B(\DP_OP_13J3_123_8774/n734 ), .C(
        \DP_OP_13J3_123_8774/n500 ), .CIX(\DP_OP_13J3_123_8774/n501 ), .D(
        \DP_OP_13J3_123_8774/n757 ), .CO(\DP_OP_13J3_123_8774/n492 ), .COX(
        \DP_OP_13J3_123_8774/n491 ), .S(\DP_OP_13J3_123_8774/n493 ) );
  CMPE42D1 U1197 ( .A(\DP_OP_13J3_123_8774/n520 ), .B(
        \DP_OP_13J3_123_8774/n806 ), .C(\DP_OP_13J3_123_8774/n524 ), .CIX(
        \DP_OP_13J3_123_8774/n525 ), .D(\DP_OP_13J3_123_8774/n829 ), .CO(
        \DP_OP_13J3_123_8774/n516 ), .COX(\DP_OP_13J3_123_8774/n515 ), .S(
        \DP_OP_13J3_123_8774/n517 ) );
  CMPE42D1 U1198 ( .A(\DP_OP_13J3_123_8774/n780 ), .B(
        \DP_OP_13J3_123_8774/n493 ), .C(\DP_OP_13J3_123_8774/n497 ), .CIX(
        \DP_OP_13J3_123_8774/n498 ), .D(\DP_OP_13J3_123_8774/n803 ), .CO(
        \DP_OP_13J3_123_8774/n489 ), .COX(\DP_OP_13J3_123_8774/n488 ), .S(
        \DP_OP_13J3_123_8774/n490 ) );
  CMPE42D1 U1199 ( .A(\DP_OP_13J3_123_8774/n535 ), .B(
        \DP_OP_13J3_123_8774/n854 ), .C(\DP_OP_13J3_123_8774/n539 ), .CIX(
        \DP_OP_13J3_123_8774/n540 ), .D(\DP_OP_13J3_123_8774/n877 ), .CO(
        \DP_OP_13J3_123_8774/n531 ), .COX(\DP_OP_13J3_123_8774/n530 ), .S(
        \DP_OP_13J3_123_8774/n532 ) );
  CMPE42D1 U1200 ( .A(\DP_OP_13J3_123_8774/n544 ), .B(
        \DP_OP_13J3_123_8774/n855 ), .C(\DP_OP_13J3_123_8774/n549 ), .CIX(
        \DP_OP_13J3_123_8774/n550 ), .D(\DP_OP_13J3_123_8774/n878 ), .CO(
        \DP_OP_13J3_123_8774/n540 ), .COX(\DP_OP_13J3_123_8774/n539 ), .S(
        \DP_OP_13J3_123_8774/n541 ) );
  CMPE42D1 U1201 ( .A(\DP_OP_13J3_123_8774/n554 ), .B(
        \DP_OP_13J3_123_8774/n856 ), .C(\DP_OP_13J3_123_8774/n559 ), .CIX(
        \DP_OP_13J3_123_8774/n560 ), .D(\DP_OP_13J3_123_8774/n879 ), .CO(
        \DP_OP_13J3_123_8774/n550 ), .COX(\DP_OP_13J3_123_8774/n549 ), .S(
        \DP_OP_13J3_123_8774/n551 ) );
  CMPE42D1 U1202 ( .A(\DP_OP_13J3_123_8774/n582 ), .B(
        \DP_OP_13J3_123_8774/n859 ), .C(\DP_OP_13J3_123_8774/n585 ), .CIX(
        \DP_OP_13J3_123_8774/n586 ), .D(\DP_OP_13J3_123_8774/n882 ), .CO(
        \DP_OP_13J3_123_8774/n578 ), .COX(\DP_OP_13J3_123_8774/n577 ), .S(
        \DP_OP_13J3_123_8774/n579 ) );
  CMPE42D1 U1203 ( .A(\DP_OP_13J3_123_8774/n618 ), .B(
        \DP_OP_13J3_123_8774/n864 ), .C(\DP_OP_13J3_123_8774/n619 ), .CIX(
        \DP_OP_13J3_123_8774/n620 ), .D(\DP_OP_13J3_123_8774/n887 ), .CO(
        \DP_OP_13J3_123_8774/n615 ), .COX(\DP_OP_13J3_123_8774/n614 ), .S(
        \DP_OP_13J3_123_8774/n616 ) );
  CMPE42D1 U1204 ( .A(\DP_OP_13J3_123_8774/n623 ), .B(
        \DP_OP_13J3_123_8774/n865 ), .C(\DP_OP_13J3_123_8774/n624 ), .CIX(
        \DP_OP_13J3_123_8774/n625 ), .D(\DP_OP_13J3_123_8774/n888 ), .CO(
        \DP_OP_13J3_123_8774/n620 ), .COX(\DP_OP_13J3_123_8774/n619 ), .S(
        \DP_OP_13J3_123_8774/n621 ) );
  CMPE42D1 U1205 ( .A(\DP_OP_13J3_123_8774/n590 ), .B(
        \DP_OP_13J3_123_8774/n860 ), .C(\DP_OP_13J3_123_8774/n593 ), .CIX(
        \DP_OP_13J3_123_8774/n594 ), .D(\DP_OP_13J3_123_8774/n883 ), .CO(
        \DP_OP_13J3_123_8774/n586 ), .COX(\DP_OP_13J3_123_8774/n585 ), .S(
        \DP_OP_13J3_123_8774/n587 ) );
  CMPE42D1 U1206 ( .A(\DP_OP_13J3_123_8774/n517 ), .B(
        \DP_OP_13J3_123_8774/n852 ), .C(\DP_OP_13J3_123_8774/n521 ), .CIX(
        \DP_OP_13J3_123_8774/n522 ), .D(\DP_OP_13J3_123_8774/n875 ), .CO(
        \DP_OP_13J3_123_8774/n513 ), .COX(\DP_OP_13J3_123_8774/n512 ), .S(
        \DP_OP_13J3_123_8774/n514 ) );
  CMPE42D1 U1207 ( .A(\DP_OP_13J3_123_8774/n564 ), .B(
        \DP_OP_13J3_123_8774/n857 ), .C(\DP_OP_13J3_123_8774/n569 ), .CIX(
        \DP_OP_13J3_123_8774/n570 ), .D(\DP_OP_13J3_123_8774/n880 ), .CO(
        \DP_OP_13J3_123_8774/n560 ), .COX(\DP_OP_13J3_123_8774/n559 ), .S(
        \DP_OP_13J3_123_8774/n561 ) );
  CMPE42D1 U1208 ( .A(\DP_OP_13J3_123_8774/n611 ), .B(
        \DP_OP_13J3_123_8774/n863 ), .C(\DP_OP_13J3_123_8774/n614 ), .CIX(
        \DP_OP_13J3_123_8774/n615 ), .D(\DP_OP_13J3_123_8774/n886 ), .CO(
        \DP_OP_13J3_123_8774/n608 ), .COX(\DP_OP_13J3_123_8774/n607 ), .S(
        \DP_OP_13J3_123_8774/n609 ) );
  CMPE42D1 U1209 ( .A(\DP_OP_13J3_123_8774/n574 ), .B(
        \DP_OP_13J3_123_8774/n858 ), .C(\DP_OP_13J3_123_8774/n577 ), .CIX(
        \DP_OP_13J3_123_8774/n578 ), .D(\DP_OP_13J3_123_8774/n881 ), .CO(
        \DP_OP_13J3_123_8774/n570 ), .COX(\DP_OP_13J3_123_8774/n569 ), .S(
        \DP_OP_13J3_123_8774/n571 ) );
  CMPE42D1 U1210 ( .A(\DP_OP_13J3_123_8774/n526 ), .B(
        \DP_OP_13J3_123_8774/n853 ), .C(\DP_OP_13J3_123_8774/n530 ), .CIX(
        \DP_OP_13J3_123_8774/n531 ), .D(\DP_OP_13J3_123_8774/n876 ), .CO(
        \DP_OP_13J3_123_8774/n522 ), .COX(\DP_OP_13J3_123_8774/n521 ), .S(
        \DP_OP_13J3_123_8774/n523 ) );
  CMPE42D1 U1211 ( .A(\DP_OP_13J3_123_8774/n604 ), .B(
        \DP_OP_13J3_123_8774/n862 ), .C(\DP_OP_13J3_123_8774/n607 ), .CIX(
        \DP_OP_13J3_123_8774/n608 ), .D(\DP_OP_13J3_123_8774/n885 ), .CO(
        \DP_OP_13J3_123_8774/n601 ), .COX(\DP_OP_13J3_123_8774/n600 ), .S(
        \DP_OP_13J3_123_8774/n602 ) );
  CMPE42D1 U1212 ( .A(\DP_OP_13J3_123_8774/n597 ), .B(
        \DP_OP_13J3_123_8774/n861 ), .C(\DP_OP_13J3_123_8774/n600 ), .CIX(
        \DP_OP_13J3_123_8774/n601 ), .D(\DP_OP_13J3_123_8774/n884 ), .CO(
        \DP_OP_13J3_123_8774/n594 ), .COX(\DP_OP_13J3_123_8774/n593 ), .S(
        \DP_OP_13J3_123_8774/n595 ) );
  CMPE42D1 U1213 ( .A(\DP_OP_13J3_123_8774/n508 ), .B(
        \DP_OP_13J3_123_8774/n851 ), .C(\DP_OP_13J3_123_8774/n512 ), .CIX(
        \DP_OP_13J3_123_8774/n513 ), .D(\DP_OP_13J3_123_8774/n874 ), .CO(
        \DP_OP_13J3_123_8774/n504 ), .COX(\DP_OP_13J3_123_8774/n503 ), .S(
        \DP_OP_13J3_123_8774/n505 ) );
  CMPE42D1 U1214 ( .A(\DP_OP_13J3_123_8774/n592 ), .B(
        \DP_OP_13J3_123_8774/n814 ), .C(\DP_OP_13J3_123_8774/n598 ), .CIX(
        \DP_OP_13J3_123_8774/n596 ), .D(\DP_OP_13J3_123_8774/n837 ), .CO(
        \DP_OP_13J3_123_8774/n589 ), .COX(\DP_OP_13J3_123_8774/n588 ), .S(
        \DP_OP_13J3_123_8774/n590 ) );
  CMPE42D1 U1215 ( .A(\DP_OP_13J3_123_8774/n739 ), .B(
        \DP_OP_13J3_123_8774/n762 ), .C(\DP_OP_13J3_123_8774/n547 ), .CIX(
        \DP_OP_13J3_123_8774/n545 ), .D(\DP_OP_13J3_123_8774/n785 ), .CO(
        \DP_OP_13J3_123_8774/n537 ), .COX(\DP_OP_13J3_123_8774/n536 ), .S(
        \DP_OP_13J3_123_8774/n538 ) );
  CMPE42D1 U1216 ( .A(\DP_OP_13J3_123_8774/n628 ), .B(
        \DP_OP_13J3_123_8774/n866 ), .C(\DP_OP_13J3_123_8774/n631 ), .CIX(
        \DP_OP_13J3_123_8774/n629 ), .D(\DP_OP_13J3_123_8774/n889 ), .CO(
        \DP_OP_13J3_123_8774/n625 ), .COX(\DP_OP_13J3_123_8774/n624 ), .S(
        \DP_OP_13J3_123_8774/n626 ) );
  CMPE42D1 U1217 ( .A(\DP_OP_13J3_123_8774/n407 ), .B(
        \DP_OP_13J3_123_8774/n411 ), .C(\DP_OP_13J3_123_8774/n746 ), .CIX(
        \DP_OP_13J3_123_8774/n769 ), .D(\DP_OP_13J3_123_8774/n408 ), .CO(
        \DP_OP_13J3_123_8774/n405 ), .COX(\DP_OP_13J3_123_8774/n404 ), .S(
        \DP_OP_13J3_123_8774/n406 ) );
endmodule
